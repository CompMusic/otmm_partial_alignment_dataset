BZh91AY&SY[�% i_�Px��g������`�X�׵�� #S�����l�$�44#@�?M&�i��M4b ��J���� &0  �&MLL`��f�D�����2   � �Ah����B~��  ����A�FH�6�ɠ ���-��q"%�D/@	 G��I킐1��Q�P���;(
���(pf 	�Yg7����cɿ���i����swMwk��w7wmw��9��_1�-7�]�z!��`�:���e�W��\��,XwP��S��mS)�A#�Y,�2)Rfc�,R�.\��3��|{�.v����X�N&,�l�k�ᚢLu�S����-���u\�#
,�a��,z.FwV����UDKr�J(����ًC��ك��d�ٰ��r�8(ɚ�<p�
��`E�.+ykWFw�Q�"%�6u�w99[v�薦���V�3r�$���CЙ�4 )@ eG�D[�G�6p�3�j�<@��qB��޹�cS���O�p9�)��Y�V�r)�z��)�� FGVQ��V(8���0��d&$��c�� i%U=�%��3��|/l/��WP�La���%�֙�:��`CC�8��T����?4|d��S��Ӳ�Ri5��]��H�`q:��L���&9���R�7�#_`���ڼ��It$L��vą�-sƅ�W��T��q4���I�O<��1U;;u��z�\GF>b�K�Oo�l9x\Q�Ro���8�c[8,��WQ���&���ة��K8��ˇ:>�21�	;�����fZ\P!&aE�b�hp�m(��<�ZuC[߂�m1�Skإꨔ-3!ĥ��p8~JA�#X0n��}��3A�m��!2;�@HR����k�woCq�������b�ݿ҇��v2U�t�#�O��1:\3��H!�u���5xF3�N*��m�u�h(Y�B���Ҥ8] Skp��`&w$����ѱ)!� Cm2!q����A�o�)�?�D�ii��M����#OY2aG�ph$0�q��1'd�@؊��t�:��jZ��@j(�[
*�H-lbX:d;���W����w�:�6M�5�#ƏTyݼ��/�f<ʇ�}u���s�[�t�(R�G:�\|5~�%EcU;�c���ih�[�2��1�DHVkj��1�u�ok%���ܗ��G�'��~��`����ݍ�>$�B]f���(���H8M��5r<oS�`Qɬ�v�X�&��8�$Y]z.�*\3�u����g��W�t(AUA4��*�ąa�F�'}��B�����%����`�4�&0li��u`��A`i�;�2�"��M-
}�<IS)AF�FL�}F��^����5�@5��ʹl�\���H\H]��J��8:����zl`�B�=d����1L�ԶGe�#t@�
�i�8��E�b����Mۉ͋c91U��49���J��HV�I	������P7}�8j���,��jgq�-d���B�ܺ dl�ġ-nEIBB�)�FEi�KCI-��[Rf��lR�@M��B���^�*�<ĸ��Bl� ��]9VfT˲�ꋪ'Yf�Q!2fT�w��	�ҍbB�y2�m-HI�?�]\��K��ej�A�hwk��p�!�����tY*7� b����q
�4=�"���r�Y6���E�D���@9����nc��\�L�K�~�}5:Uh4F2�P��T��J�wxX�LJ�������9�f$���
��g�L���\*=�t1���iwf��S�r��4�*38n�m���mU�/��5��C9#�P����J��ܑN$��F�