BZh91AY&SY�c�� 
_�Px��g������`	^X�׾�ʪ  ���]��4�{;��&F�OS�2y��4ڍ!���L�D�#M4��!�b0��7�$� ڀh � h  ����E��=M��@�ɦ�FCA�Hġ�ɦ��I�2h ���=M �#EM�)<��@�=C@  
��Ң�(�.T
 M�E�V���V4���o�P. �A�`fN�S,m9�U���1�v��g9�{�����333�������wwwouk�����r��p�r����4��50"�q&NL�J2��F!%A=�qڐX3iMdR�k8��.<��i���/������s�kP�`�fl��0����\�r��n<6�/��2ٛ�V�4�jڊ��-K��[\��2]h"��Y���uߢ��1��V����y�G�(�3��RBG!M�(

��ŀ�7}�����
�0�|ϵ߶�����u����z�-��S�v�\51xbb𡒬˾-ta4!k&%F�Q���߶38��Y���"�����c=�`P_�4>f��K���=�71��\[ux�����q�;Hk�|!�����"6s�9��E���`��T��6qQ=5@R�u�۲�jm�g:p;9ۼ(�]<�#X*���Ex���#�r��[�'ޱ�9 F�N��y��t���q�p������@r���\D&s%��MǺ�0�	W5m�*C*�;��{Ƥ��q���(&qK�8@� >�:��#�S�)z�b�x�#��μ�D���ԛ�k\8؉���Rut'��i�9K������F��u��L܍�q'+@ښ���y�H�xmxP�i�����y'���<>�*d���+)�xخ!s]}z�K�Z��K�ݐ���p�h.�@�'�AË�V go�蚫i�r���Us�G%�õ9���D%��Q�v�����v|x�ހ{RU�9�������he���=5�������Qț83p;ƌ�S�t
����=�evz���^���~�H���nN>E���9�pOJ�Oq�D�v����R��l�#_�����/�g��t	�3̻��o����ߏ�+Ԫ�4$�ݧ:��G�D�椄�I8��r\<(A�)��G�	J�77*�T�	r�ҭM��-

�6"#M\��+C�FX�eZ�5�k*�жBQ���N6�"Е��W�[樗�D�.�*�d �&��DW������Y���:U��}�h�1�;Qo����e�{�N�O�橬l�x�~��MC��ٴ�k�vH��R	.���7��Ќ��S����{��%J4`���� ��7�f�g!�\T�(IA/��C�߬�#�
�^p9�ӥ��٣�B���5R�\C���W�k�!V!d�����f�~����&���TԤ	,��I{I�hE�F�]�)�d�H�$� H��**����+(��ٲ]��W�`�=�<���K���C�,�s&ZT,ˠ��Q�p�gv��T����K�_��5ގǭ�[���V��DV�#�8�;�F1�U.Mj#nꠕJ�C������~7�RUʶ�#q"E������`N��&��J����a������a���>�\�k�h@�*Cf�W߭�N��(9�ZޛC Wq�qp2)����+�Je#
a#a�D���A�ix(,㝥J�p��*8)JI^�5����c������֘�9LAXR&ͷ4fL��%P���3 �?�x����ej��3�e,����p\��`s'BJ|��+'��F�Is�%{~�n�:�|�۲֋6�uI��;A38�9Nn͐[U,^k��Z�[����ϣS8vG9`34�z��֧g`�(n.;\�`cl�,LX$��^
��}��g�ynbhI��P��b��m�d�=U�tW-��h�i�rD�hm����S)_���!h����"�(Hs1�]�