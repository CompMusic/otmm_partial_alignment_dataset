BZh91AY&SY��B w_�Py���g������`�{s;�� ��IҨD�2�2d� �i���F�h���L�T hh     i���ިz�4h �@  &�&���
C�C#�0d ڀ� �`�2��E�CDj~�y55=꧔�OF� ��~�=M5c�$Q��B@�����e"�$���)���� �0��*pfI
.�&\������ӫ^��ݻ�@� M�!��oԻ�7�c;�R��dv�j��!n�M�B�@ab��m 27P֨�w�׶d�]�紋�x���F��NT�?y5I�V��6�LH�[e�$0�9�{֯<zF�X�)���������1j����+�?���zތ��ET*c*��$J��!���hߠ��O�|��c~L��gҚO�Qq�CWb)��}���U�D8y"X	H!��"]#1*R�(��#������`�5C�"�gX�8����\#��l�;)������&��(y�o`�����$�pE�+s�%hUN/d�x��x���c�c�ݰ�\�nvWr�<A�f+3|{���'ړ�X�F�rf�dZp��� 6(p=	��9m ^��n<�rt�0�A'R��l���F��Q�v��
���,K˵�騜�/���!�TG�\q�[➓�M��iّ+�E��f����;�ە��Q�3�r�8�Vq����~���Ae��ѡ��(c�7�`�1)�8�f��Y��ə�l�rЭ�i��P��5��ws&-w�$�DO��|��E�X��;Z��n�D$8q�{j��ƎU����Y7�'��w�^��7n�7N��:
��@�+j&Ｎ�xfqp&�A�
"���A���jH��f���VҊRf���I<n�Tt]j�ܳ�&�a�
;��7�l0��2]�@c�-�.���p��SmK�f˪V� ��M�g{l/�i�3���Y )�8=�&�_�ـ\���Vׁ�T�F��փ�)i�vG6rPeg���
)|���!�q�N�{�Ï�F41�H⛹[м�:�s�g����|�b]I�4�wY(�� HU�v�=�~����x1E�O�SV��H7�A���;�'�ɄS�xo����" �������KG�>r� �gcMK����C��"M@�(�	�{�U:�!��<Sٞ���ޖ`P4�
H*��4�X�D�;)&�� �=��MAZ񥲔�4�.��F�ȧ0LA�������2�U�cX@�6 �XLp���B���{P�7�[�q_���c�Y(*W�HX�n������x6"Jv\c^��.j�S.��Y9VVғ��0o��-�k8�!����X�����B�]9��i˙_��*�|O���&�'QzL�m�gBdO3k��Q	�����H����&&6	(k�a�	
�7�(%[���MR ����&�%��LwsLG7���AX/1��co2lE>��yd=�l,'`��_	�Wk8�܃������@� l�A�(n!�G��dT�����z)�U������Ϝ���w�;.u&h����^��uq��uVj��-�L�l��`Bɸ�Y�mnf�f4i�z)��j4ڳ1l���v)���lɲ��|�)�m�"�k��V�OF;
69�R)�ű��MtM����j a�ыk��1?�� �{�q���}�9��w$S�	o�T 