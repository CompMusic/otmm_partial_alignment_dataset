BZh91AY&SYs�5P B_�Px���g������`	�����   �ⵥJT$��艦��4i�6��I�F��h4 �EF m 0 OSʩ�`FLɀL �d�� 	OI	Hh 44    44d���`F�b0L�`�"4���O����S�O)�h ?T�%���� DTh$ ߞ�ף&��hu@P��'��b��R����s�r{�pǷ�;��gvU�c33333fNf6e������̶������i��+��]�a.�ޓ�&�d.e�\����2�R�eI��#^�1	t n0q�&�(o�,,ė���H3��EN�80g7/X@�3�2���)K�<�X�15$I|���,�X� ���<����Šk.rt��c�@�
��ء#"�_��apҰT?e$d38�T��V)N0��"hy�T�y3�@fA*L�3/�� 4���r��[�
��jǅo�y�tY ��+3��RǄ�.(R�19ͨ�(�3�5jӶ�4 0H� ����π0#�z���y�cq1$8J��ˈQ��rR��P�.�jۛ��lk��=J�hȣE�&� A�JA=��@K� IJV�fڹF!/T�8�0Tp�*R�N�@���8��$D�REQh���^s*6��hU�T�&�pQ��a%�R�X&lR����MZ�SC���ę���ė(fH,��
T,@V�f�D)�<m-,�T&�(�לd���J��1�fR����f۔�
�C�X��6� 7�M�<��Q������w4<	�O����wo�����Ed�$u��!)�����ar-�{�	��	la8���3U ��O4�n�7%�7(��.,zl����7Zz	�<{n*�A]]Jڙ���
���F0�x�U�#AE�~h�;�J�u�4C�!CFxE�W��H�,�!D�E����ax�ܕ���M��mС\�����Sm�jfm�I�$Wz� n
ʮ���9�}��^=7�8qu��t���-&��uYd���dw�D!@e�q+�1+�#u��&G%ﮢ��8hh؊��Bֻ�����rSB�L�������mD��GE��o��Ct"����E媪	@���W��F���c�y�P.���}҂�Ւ�v����U�(�d��I�F��A��kD�U��8�4��@ĖH��c)�37��ECddb2H��Fa���$W2�i�n��(gmJ�k4i�4dCMn�k�����X���	6N����Y<�m�'�D��/�����Ch�N��S�U��|p��r�!�M����uY�vk��V��kR�ҭr��j�۴���`�|(�^B �70I6�y 8�I�Y��ۢa�N��@���^����3Y״\��@�峄�O��ѱ��%�\�qA
K�mA�;�]\��&��,S� .6�-}�V0����}9��`���`�j��Cb@Z�ʨ�TТ�X�E� s��FNq<��du�g*2Q@�!Ӹ��
�~���.\�)U 0=��6a���{,	��\B5[������jd��$�<����kܩ1����������nH��ݣ���q�E�Ɏc0�8]��lʫz 3�� <��|��˲����7�-�jh9q@�ڼ@hىmѮE���-̀y��E��KK�#P� �%��`A)4$͌���ƚ�������LpDC���!�+�ԙ�2�Ag}���vɛ] ɵqú�������h?Lt��H	0����u�u3��-�<�]�6A����0�่F\9KJ�{D&1oy#z 2	 g�гun)�:��f�VtX�m�&c� �I��b5{y ��0h4��ճ�U
�Z1��2w�(A;[�� ��|AJ���A�����s�S4��T�@K]�&�|��#G������O���V2��Ǻ��!p�+qG0O�����e֌k��Α�h>v�Q�WC�.�p� ��j�