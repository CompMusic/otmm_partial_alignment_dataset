BZh91AY&SYl)� 6_�Py���g������`,�ug  �Ɉ�0�I��dɡ=F�����mF�h4ښz�4	(COQ�C@    �& �4d40	�10����M2��   �& �4d40	�10�"e4�4)�Ї�4  A�@I!-�!$�H�4#�b�������M��L_x}A�4����<���I)\�v[.�����KZ�&i��~���e݋�����\�jeW��Q�YZ���P��c%*��Sˇ{�-B�>�ђ�&�I��"^aDIr����;'3�~6sf���vW�ơX"�T�K"�HPħ(lAsq+����ɭx��ML؞$*�r�.CqnO3�i�}*�v� �����L��좰�	2E�r�۶l�e&L�e���C�x���eO�;�nG])��$tn�Q#��x��1&h���t�HD�q#m����c0(,<�"ݪE0�^UR%��`1���P9nmf,����MM�����KN-� ��,���� �`g�F#��h��(F����F�$(H\*A)p��I E-��:����4t��VbV؟(f'l7fc��3��� k�6&�gB��K�a��>��s��6�7��D��,�ա�ejB�+�{g�FIՇY��d<�K�,>A�0Ǒ�w��2�Dc�i��T���*w�w�8Ȩ�+ya��/f������HM����Fuհ�OЌz�eƶY'���b���[x��4%ԍ�J��lr[�J��Y�+Zs�N1��(("�XV��r�J�ջ3s��R��V���J���w|�	%p��|y������E	>gK���J�4e6��Ðw�E
tN�S��Q���F*����Qw�dހ�ە̧'83��u;�hыe�|ki&��"s%h_�؎?
oB�b$r���P�1���`��9����0�ݓ7�k���s�����t�QW��4P��x�ɯz���d�T�ndxڈ��Z!��Mk���
���ݩ�e�H�NG[��K�!"��r�UZE(QXʡihka�����
���˿�
˶�D��p�5AL�f'h��[��<��檎��{��>��<��w�NO��+O��1x
u1t����Y8��6==����`�wY�\Y2��5,�>R��� K5�L�&�o�[	y�K����%�����6v�h	t�M�|��Q+�B|㊙�����Ɖ8�7��YK���P[B+[U� ��6����u���7�U�Q��(ХR�)H�-!ԄUDZ,�R.M!F]8��
��9I�0k�i�	@��2T��v���1���W0�3.��
�Dz��Ǆ0}��!)9ȶ<��#o��#q����?.�o=��Җ��v�!K��LEu�W��|�n�+����&�6.6���M��m
�:8��f�$�p������'h��j	��@K��Z���JY��@����.��u�s,,hIj6�L�a!MP wHpD�K�	�!�t��!�������p @Db �5������H#�>3$������b���(��/�p�A���H�5=��P�+z ���#@	`(@��%�>��2�k��Q��."@�����8}0qч[k��M���Y4iĖ��J�� %Fy�e�8���0��ҁ �㤶u*�K��l���h�>����Fh�'������3-*�(؁(81�t�+��]�f�k�6��G4�j8o���"�(H�� 