BZh91AY&SY���J �_�Px���g������`�z�:��HH��ڎ�F��BH� �i��{D�hi��=@h�=&�cE%#M b� i�d 4�A	h  F�   $҅F��M �  M�101��&$HD=x�i)�~�� d����	+���$"i!"�H0H ��B�L�U2�����  l���b �@]�]{߯�����s���WL)I$�wb����%���5�C��1t�Ai� �2ﴗ��jd\��<�J��â�����Ѣ�p��3[���|��).LK��s���8�����7t�mHP����S�nX�n@��Ap͑��)2Y�g�le.s���f3Ko!�8׽&g1�Z�� � �bܸ�`V�]w)�M��]�^��'H$QJ�����J�ZuD:�Jc(�{�dɆm]�umN�M{�,�-Ϣ���s-�B\@F@�,�Hd9����8qJ!'.���@�$f,��iJ�GN�����t���D	�א�>�]��fp@Rژ9 ���rbN7_�z���������d�X�޷-:L62o.�%�� ���J!��s;�髈̆���B�DN���mc:����x��W���� ���`�&�"f�qOC��z4x�q�L�y/Mӛ5�j�Kb�KZ�ظoa$@�2.�Dq����PqMG2[&����� ���V6#4M�,g,D�ĵ�b"��$1u�KE�NH�`B�aUS�Hr��g�㥧U)ңA`��MX�"Y��,�S����"n�\q��9�^�R/�*�x�U�A�R��@��.��/W;^3�y�
�d;l%�-j�U�8w�I����bB�[p�jY�!i�(]:��e���t���T�.�'Eps8-��w/

,�Ak�(�j��:&��iX:*`�W�l@��XH���en��~R]���(v�����iǰ�G�� ���R�ɀ��{���z�kEt�2�����y����5s��cN�=�����k��u�E�*�	'?zo��{�]W��u@�ë��7��b�VE�p�'u5�k	���E6dnc��:�
���U�L��seQTS�X,T@X*��ujj�f)QT\g"���hz0�����G�EkW%�Є�v���N�3��q�V�w9;��_9�����/��;#͘�]��K��MP�J�D�v�y�WKF��L�(�UߟNL?-9�i����K�X#1��� 8
U�,�áZadC�4��\G��Լ,8���Ͻy/���Ƕ
/��c,�� ɠ܂�]�&�PC�U�s|�/����hR���U�	ds�[*����RE��2��۬X�0RE����3e�ڌ(rA ӮN,�2s���*b�_���Ҡ	5��@�]�]�	�3W��T��Oh��Ao��	��K�����,҃��,�pd	Cr+܍�pR��Q�3)a�;�"�ѥ#/�d�TJr$+��\lz�E���&2���nZ�n��(�e�Z��
�:�I%#�	{{W�����DCF�X#�W�4V�2H̄����22M�VN����i k:�5�}��cEP��`imT	=�`���&��r&�S]��]M:ɛ�� �&��l	�捀%۸��=�IA������_��2�mA����Z6\��l�H�5��Sù�c��7��� ��̦�.z���Ԋ6�qI�z�uq��j�� �S0rb4�ڶ|d�.�D���)qi�S�A;S�p��K��²5'
�g5	��a=g	AIl���R�]�H���x��^)����샪��阛YB���R�o��}��7*Y��ƿH�3�>J�%x)�h���.�p�!	�(�