BZh91AY&SY�;� �߀Px��g������`�:|�� 0�3ح!�M�zh'�4�i=�ڌ�I�� �S�EP�@ � h  bM   �   $҄(�=F@��F��@b���昙2h�`��` ���D�M�1�oT�H4= �M  �z��h����TI�)b(\� ���I�&R*��	P������ �*� "��[>��g�yÏg+N�w�u�R�cb������U
�����[���$3*O�fLt�X�����*������T�E��u)�v������j�e��RpB.S-%fR\��-r�-ɜz�ɞ�/��\���7<6k[��!� �'����Spܰ%��J)��rT9A%�čn"c'�|XQ $VZ��B5�ˁ�F����t�֯1��f�D�"	R�ʩ��J�Zut	��D��xz'X1���od�OK[o9��x9z�8�xx�g)	�,�4�Cz�]��"s���o fd�E
���B����"����V�0���;�m$����g��!Q� q4F�i�K/Pg#�W�A~$��'9�0F�p�[����*�af�($�)8��6��ޤg!��˫��C�Gd�@��#E�[+#�UUgT4
�;~
�"�"/\ѶnB�d-����MtZh<ƶ��e:[��[�m��u�3������!��Ր΀���Fi�j�*s�l�ع$L�U��d5�GVJ�!ΐE
��=s3�2��e��bAM�%!�1�Ba������^�N3�QOj�}"`E�����lLjZ�91�B�:-jYa���AX�-ggԇ��/��.*�`r�D��ڊ��i$1G�ټtlPB�`���"Q���fDLw�H�_N�=���o*����.T�K�+_=>t���3ʅQ;��\>8��B��fʵ�:�YQ�*9��jR"�//�Ŵ�U��3Wh2@�v<�����뽖�uz�����Pzf��[XV./���է�Pc�^���H+��T���r�9�L�^���vE�̭��n}��۸�QW�UT4N�k�9Xï�]W�ƃ:�I�����>d��ꩤ0��q&][XN*Y�QS���n�.��lAE�e*˦WE����
)��,*0ᕂ�*�m�E��p����إ������gn�<�hC�|��Aa��-���*�7����8�rD�{�V߇��X�g�N7S��~�?ۮl���*�~�k���.�c�?.�ӪRmA}��m�[���_�ց�b�e����+i��4[4�@�$� |��K����5�9AfÏڽ�������ʢ,�.�hpit�K^�A'�˟��4��c���J�-�� ]~&QIq�������Ξy˔L���[$��T)"�@FD`�YUL����7t�3�������12�J�$����,���Md��Ev��m��6ñ �s	�	~�B)��u,���V� ��6�w�#�r����5���Nƕuϰ���3�M���w��|�$�4�Pr�,����s��l�ųG�XG�]5�}��o$���*���/���o�d@���n��󸫴h�#"��%y���"���U��i di�	,�$"j�	c�"`%�)���
���'	��C��j]��6�D�s=�NF{Sp����������x��ܞ1���C��)FW�=A���*6�ϸ�82An�т�މ��+f{=}w�znn6��M�D6X�dN���+��{�?���ꛡ�Y�����]�R����E�mk.�D��ƲRD��аH/���s�;X������PV�ф��b�_HӺ_�r�XuO&�CXġ^�Ab����ݔ����M抖f��k������U?��H�
g}� 