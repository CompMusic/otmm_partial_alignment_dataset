BZh91AY&SY�҅� �߀Px���g������`{��` �.�iщ�R��	�i�I�a� hi�Mh�4h$� 4�@     挘� ���F	� �i�T� �  dd@z�#U#FMA�i�dd�L�hh��)�OSFM��4  2 ���.��H� �$�O��G��(H�I~��Z~��H
r�� �Qe=^�oQO������?&fFfffff�����\������9��wszW5U��㑰�'/��S*���+�X�3?:u�\�:igcU���$�]��d���㸻QŦ/":�Lg}:,��v�ys8>/{	#CW?Ȉ��� D� $��]��;��T�vܫ��	�����R�)��$��N���0Z���2I&L�eU�S���I�]��FR(�������v�:cNE�si����w7w1��D�j�K�o�fpa�-�.뚙LwڷwQn�[32��_N� ��dS%ߘ}CIV�`C�c�*�&���@i]"M`�)�ڦ�m��0b��ZӰ��"�è�!8B#�M�B�(�@�˛X$����;�sZ�
�D������YV��e9����G�M�Z���+��<�Aq�Y�W��%D�5Br�q�kc�8��{�]��E��7(,�E�����wb�N���j ;�Q��A�mO8�+���K��P���/��Gn�qf�\w!�� 7�v�dA�2���EN��t�%�0�)���R����rw���c�����E��tATl���S�1�D��4&�,�
����E��(@j�J�p�[n��ij��B9~:^HXWyiSdA����gp���IQk��]o3�mDDGn����H��v��e�p5�`�!%z��*�Y1�S�:
�tn���KM�A�j�QRn���2�4۱T�"�qO��x��� ��sh9.��f5A���8���m�  �N>^�'����ӃY$�W�q\U#.ܐ��좑`<t01���)C�N�]a�T�TQDFqi���^)V
	�f[� �͵p�iF����֗�*`[Z㓢w;ޤ�n��j�-x��` �{�1�{�<WY�]nXx����u��v�?���Μ�^U���Q͡���u�m}3�F@q��Y 5��M
�n��?%������&���r��sg����:��RI*����-7m]+bI.��ϕ�؛�T_M*�\��(R���*c���|c����ZܫT�X��lMXL��Lr4��bF�p00�##`+"E��@���1� ���(ʇ>�|��I%�ڄ�	���������y�ٌ8
���I/��#^�D0�O�g%v4�=�E�2܎�5Bc�cNB�c_�x[:��o�Y#�iV���q��-sվ�Vi$�X0 0ت�`6�#�p�E+=�F�˙$ ���Ix���"P��N �-I%�nY�Z%�� /��&�j	%�!�I�f�EU��#�{pD$(b��Y�D�	�f=��n����ɲI@�u��$�x�GNzM) 9��џs%�ox���yb;��lR����P mA����I%�Q$�jyy�4�aww	W�.8���A��p�p��3�8�C:�ͷ�mV�,c���n�lI%e��w���%o�pv�BCL��KKZI.�H�l�ѫ��e�x�� ��C�&E�$��JI � jq�
���_Yu�����<�� s����.�p�!3�