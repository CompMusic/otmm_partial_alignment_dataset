BZh91AY&SY�#�� �_�Py��g������`~����  �\N+v��I&�MM��M5<��S&C�3P�m&�����@	$�M       9�14L�2da0M4����$Ԅ$�H44zA��4   �T�����G���h� z�  H���6�����4�@  �"�]x�"*R�b�U��i�e����!"O�9��x C�%K�0�0;�e�a~z�_'�u�j�U���U�����UL��e�9������mS�4�<0l���̻
�Ǟ�5�M[�����J�fjʹ�O ӄ�R�# �B)D:�fB��Lvy�Y�d�fL���#�������"_v��()���`Y�����m(��
&���HI���P�A#����Z�],-�׌4�P��ĈM�mOIo9R��#G)8����0�SM�$Ɇ��?�l�1�{Gc>�($xw̶4�����:���%��J�Vp��8b�A.��f��<]FJ�
���&�Q��CA1�ޚ*�3tal���f�\@1�f�!f�nq��&S��u��N�q`������r@|�*��,P�东^���1 ]�:з�J:�[���PBi
%]�j�$�
���[��^�.@��s����f�l>b�����pA��U��`�T�.�)E(:)C^B�9(U�iUYq��{8���rie�2D����H��[��ٰ��&H@�u�E>M���Z8v��.��YF���f��ѡM:.���3|�r�f%��KE��:9A�Z�N#m�TH�9��9ܙM��$v�;r� 
���;2��Ã8l긡5FJ!=˙�#��-��'�ws3w�QϢ����+VN�JG:Iਮ��.6i�.������z�ƌ��wHN�6©��EX`���J�ӹ����%6-�D����#��D1^���lXz��".;�0��i�=�eu1p��j~�iYɹ�Wh2�t(�j�v�3��h�b����7�},����O �����]qE��]��\\�h��T�SȸW~2��*����I
��HЛ�=ӓ�dt,a�1.������h�MҪ�^j�B��:Yj�b�b+�(l)�B���oT�Ɂ��.���*�		�T4e"6Je�QP3΃��4��xa�0��ݛ���H�����s�^'.SL�6��׬�wl�`��I�<�ς{X���'��{h��g������/r���	_[��>u翬^2[�А�hń!����+M�Ϩ��M��QG)s���Y��^q��q�<F��~�	�0s6K��.��L�����w��$R��ZL�BM���k˂��-`߼Ud�YE�DA`�,�AV�*��p$ e�Td�^����F��:a����,�zeiNb�3`�l��4�"��w5D�1��xI2P�:�!�=#Y�rf�7������q��[��>��9#��E���7���pl�y�0�BL6S���ݘ�s��p�����Ȯ�I$��B[t�H��8�'CU#���B]fՖ���#��d��Lpb�z�L9[^0p���M���f:��T�I져�̴��L�&Rn�0�d&P��P#2Bj�}2�[ts�/g7bI'`��upƾ�2�\�H������8�G0�C.��!*�	q2/��Fb��N��%�fꉶ�9-/	ɢ&3�pr��\ps��Q�Q��s�e�*�I:f�S���²-����,ng2$�+�:L�+a	9'��	
�w����\,�Mo`G�K�
Jk/Qo���7P^��Ε��a���1s�I#�Έ���"�(HZ��a 