BZh91AY&SY^� ߀Py��g������`>��  ��K&,���BII���I?Dъ~���F��G����y#i��S@�D�    �&�S�zh@@     iD�Iꞣ�D��G�� 2 � ���"z���h �@�h2  H�i�F����S�6�0L�@Ѡ4h�$���@H��aP(h �~���A�D�I��x~�I��"Q ��*��x����������+���fff^fb�]��M�f>]��ݵ�fV��/��m�C����uX��譼t"Ld�rjDJC�M�sQ)LD"JT�hc)M�m�"D�$��,)�c��r3G�T�ФM�|���/U
�]�RpQ"�S�0�,H�S2�2�d�!���ZځF�lq �E��� /
3����.*�ٝG��rTUm���֐�<�<s�"���e�nHG�3ŝ}]�B1��xY��n��>^�>{k�gWVt���1�u�MkL��Ш���(��q� �t(�2:!�(w�N��~�cy	��HW�Ëݵ}��2�� �K:h�l�� �)���	�L7C����Q�fHM��@�-��JI(PQ@,�ǈ����Qe����+���
�c&C2��A�!;��*X�N��e*�:�o/� e^����pC�z�zZ�L�mρ"*&�� ��R�eZi�����`:If��R�8eވ�l֗[,d	8�K��\0�k��|g�4Y��.�8�rs��޼�yvW!ב�`=,�uM�'�#-iY�vy~�iS2�r��5n�Vܮ�� �s����)@�TE<;P��fga�+�2*�3��S�'i��L����205(!^��b�E�D`�J�2¹�j�X�� >K	QY��� T�$t�M���D΀�^��67z��VI,h��.�kP"�WN�m�vF����c]@�dSvb�C:���:�-�v#ja����5�ƾ<9��U"�&�a��S��L$��,��k�[D8��x2��2t]����=��AW��!)N��5G����Ȓla���[q�f�	]�ETٕQp�¶$*J����2`w��G�a�6���Z1��+RE"0�X(�
����֓��0���t>�t@�p��z~���^C��o�]>�n݆����:�6��
Lgu^^S����Lq��;�t�ص���M���5�&5P۷2��.���G6$��C�Ma��t1��2���l��C��	:�q�
�ŴH^���[�x�sri�0�Z r�y+�*�'Og��{�޸���"�hF�*R���91į~1��v�Rߙ�I� 0PE�d �dE`��TVB��h]�SIћ�چ�6�(�"B�)�W�"g�1=�7�Ƒ�,�	��*��B�P�/�f�O�q�$�~A��t�y��S�q�N�Sf�~�y �i��ۜ�i�bD�/��
ѝ�Y�l�,�B�X�!0ؖch��X㲅��Q�ĭ*a!'�D���\�hӺk&��P6	�ִO��3���$',���˓�)�$�z�s1&f�F�+F�HO=��<q���M�Q	�E�&�+�a<	�!{WI4�t�^촔�$�-v������j�X�h�C�!�LRA�a*k*4^R�	��*w"B���2�=�l1Tˑ&��Hz�-�Y�$�ٜg"��lutd�
�pE��� �<sF��B��-��B�:,K��aז��aEF$.��/&	у, �ɤ��B�Ms��"�V$-��ZM$(iI
��n�ka�h��J�2�� Ɨu�F����.�p� �&�