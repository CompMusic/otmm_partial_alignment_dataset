BZh91AY&SY@�x� �߀Px��g������`�{q�}�HP ������KM=j($���L�cSf�M��ѓ �Ri�@      昙2h�`��` ���MD�)���@щ��a hѴ�mS@Jz�&��  �����"��L��
l��zO)���� ���9�iJ�)h(\ z�}I���@=2B2����ѢI'�2:���@)k�Əu��q�-�󮺪��ՙ������������MUUY���r7�Ꞑ`�9e�ORW��W
��D��]܇n%i�M#e8@VA�e"Ju�V��;P�=N3���;��յ��:!�v;��A�xD$x 1*A!�����+Q��W%�u
g6Y�|�jt�8��ߟ�B,]��z��x��ʢl.6߁%�	�̔n���8�TTN')A��D��e�͐��^���N�z�o�6���;�}�K2�1l2�,YAY�����/V�p]T30*)��hq��R�⺢ G;��c!ɉ�*�G�*f���
�l!�|��#r#3$\C꼘�N�A�{7P�҆0�)�ЀTJ�\���S2����S׭��$9&��P�ͧ�4��Uf���:����[Qo�<��+��M�f{�=��C=�R-�ҞHe�� ��zv��8)e
B�JB� @XQ�r��\HF`U 4�5�GT;��`�8.'qr�@_�*�<�ɒ�������35&j�+j�2��`�BI���P������n�0�\���.�e3
�gK�!��X*����/'eո_a�NT�&�[�e_t������hy��bD��p�<���?�[jE��U�v�W�;��u��N�C(d�.�j�`n�㑺-��#8���
8��,ʹ�l
�D�����ٱ%�a�8��ľs��.o��A�ܘ,�Լ��Y������aB81���+��-dх����CyM�`yc��s=UGm`��.���F�VI�1LJ��t�\kZ�p��1h8IQG��UDl͖[81�0�*_%f2�Pjk{�:O��(�+�UP@��;5�O��0���e>��T��ە�>f�4�h���M!h��T��L�P�UAFq��5�T�2�TE"�x���d)P3�M���!L��:acz��7C��ٝ��1���̵��6$��Z�Fn�l:�;�h��>�z�^o��}殌�:��#x�yh�UQ:ӳ�т�ka�c������@̤415����6o�Zɑ��ꇵw����D�D
I$<.���s� �'�6W$�f��M$,�/��Ϟ��T���ݛ84{�q�ҕ�P�\�Ua�~�	�N{1�C�����:�;S�*TN@"�ѱm��q���ۊ�Mq��t:0�h�ҭ1�`���s*���(mCC�&�-�����D�2'�y�^B�P�������1T[�魊�Hl_p߯���B�4X	ƨ��\Q3Y�.e��~[$	DȀp"��r9��e��!�D�
P�~��t�R1���P�[�2����Å�q*�}*Y��`Z�I��VƯ�`?}�{��e]Z�˔B&�,"��B������Ӥ�Z�9䱹:B�G����!2)�J� -�'��	/
`��� F֐̵@�Mxvϰ����DtUR
���2o.l��n���7��qfn�i!2MRoӥ �[ؒ�� ���^	(0��x�jv��8^� �B��x�� �(zy�l�xl��� ���=;SR�y��B����n�U���j�rC�J�6I3M�Sp�0\��fg��`B�`(Ӭ���KG˼�D	8��$�/��x�H�C��U;M$T�B�8��P���$o���� _��
�o�3*=�3�9`.Y"@%=��6���OS5S�c_'e�#�)������)�3�0