BZh91AY&SYf�r ߀Px��g������`�-�q��e� p<o��Wv8BH��=S��?�b��CF����F�O����@1�   �OM
���4 4     i&��jh  @  ډ0���&���4��    J =�M�  ����f�TP�����w��-�*U`��<��0"'<���̄�r���o�z�ϲ3��q��Ye��kZ֪��������������݋��lH����Zp*0�p�h��
y0�ItŋD.�Σ;�	�s�IF�Uh�Gz��Iڰ �h���r�Z�$�������20�J��1FRd;	\���ɺ4� H���"�}�!%�e�h�}p���8�����(�
BlV�N�~ba�@��^��#�����V0�nM��K�-�L���9�3�:��5�����H�%�*���@��j�U�tH��a$(�H�Z��r[.)ER���j(8v)���5)JQ�H_A�ūqN*H�
�E���Վ���v�Cc� A#��4�r�A�D):�MdM�a�&8}EX�v��r�@�D�z�T$��lU����p	눁&T�QLƝ-�5��ZaA �C�VU#8�V�G��n5��΅�;�"i!�WFb]���*���(���w�D	H؏��"��t"Uui�i�Lp��#d��g:��gʖ�pX`iV.��6��
r ���#g��%K�Kk-�l�A�q�y�W��=��!��j�_���\7"��u�,�W)�^$0��/��,�n�4g8շ��¸0-��9wR�s���%\dk�h7�YYRC�Ku��`5�P������aX g�7��"h�rfnd�`�8�7�;A��AJ�-X�n[�T�r�&n)��@�Q���*Ћ�8��̾@*�X���(i�k{�g�ܜyb��Ug��W,	�����N(Q�	-M�,5ذ�N�=�7_�DDGZT�:���GF{Jq�4��Du@�yټ��O,I�$4������ϖ0R�2��(2�S�YԍQ8=�� �m'8�Ȇ��ڻ&�T�K�]vT:M�HI9a @ �!�Ͻw!ڋu�t��V�d�� T	UDf�d %��PVX�	�b#pz*��D�`��g�ZW��P��J�;U@�$S7J�n��MR6�B���q&�Rx6�Z��|�����-��n���Z~�������z��΄zgX��AĖ�ߧ�mT�-Ò�����|�S��8��dp��5�I|	�W�2�v�̘}&�G� .F�$�'C3����M͂��I*Ȕ���%W���&�9���C\�e�;F_IU*P�`�l�����_͈�u�E���v{�T�yJ�b UmߵK�,���� �h�q�	$�"�2,d�H��@�SPZ]@�YK"Z�����U�UhR?��'�يe��G�+�-����ÊC@&�U�lu��Jw�w�=�
��*�X��$�)���~q�l6ǰ��bZۿf��l7k3���a��kG�u�oy;�Y�� %K���y][X���hiCx� @���U��$M���p`��(�K�oR�`��XJI�:��YXھ�e��6J��<����aH�n	��m�!�U�6�A�cG��&h��� 2vJ���`�Z �`ul^W��?�_̀���ļēŽ�O0k�QR��5N���d"aͩ4*���V���[Ǖ����7��1��H����֒�3����p�6��wY��,QY̅�)(A;R�I%2�4��Vϕ"����m*��q�_>��I'#63�{��@1��u D�%��U��$���'�qP |��ܜ�7��ݷ����6k!��Z�D�J�5���"�(H3l
9 