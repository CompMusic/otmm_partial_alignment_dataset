BZh91AY&SYB�-� O_�Py��g������`?1��p  @�U��ڡ$�OHM�����z �����M $U F�     `LM&L�LM2100	OI	!G�ԙ����=L���dc�A�ɓ&F�L�LD�OHj4�ء�4 ��bI	[��H$EP �#���WA�6�������4���s�;	���,����}�!���OWŻ��y�ffffe݋�����\����M���0j4VV�x�(~K1��LY��ý�[��!]�����u�$�*��R%�D�*���v;g]ԑ�F&,�g����"F��6�e2���NP�a����'��:V�!�e�BX��5���*W����&��+=hj	�i�H	f�AX�P6��̭Wg�xM(�oGz���1�c����ǿ~�7��SirH黼2^1�0��[�S����kP�2�Fۆ1/é.,��S!���6��G��B�dSH�=LP9nmf,���O�kS`�0$��q�zy����W$��mG]���4q0@rL��	qK�:��a	!BJ�R	l�*	 =-�!w����u�r�4�������OM����	3���#��&ä�٬�@��t*t�ľ�`��A�"G��'C�%���YS��92kh
/��3ÑCl��\<Η���:T8;&q�<�(�WFj��c�i��T���Ts������v�t~7
���^j������a���\�1��I�U�Sk�g
ۯksA�3��V� �|�8E*��ac�˱:�ZA@��gG[⒫��0�P�KB��dɠ�	H�v�N
6`����]5V�]rÄ���_T��\<�әxk��B�%:'H@NʜEF�c(iB�]�l:?8 D<r�78�gx7�Y����8b�B�f��ʆ�-ܫP�L�a�2�g(4�Z��2���G�NP-j8����k�d�){q(/�z��6�M׳�G2���A��`�}����~5���S-���j""T��6C�B�F�.�T�07jn̸Ii��uiq$$Q"�nZ�J�B��
;Il��iQJ��AV��@��M��݇�8�/�2׳.Hbl��ʏ/Ly|e�����~���}�?4��*o%2��O���N�_>��]@�F�����Tms� %���gd˯g��G.q[��@�h�B I�Tx�ti�8r�nrM� �#� �UŰL�j�[n�#���PE:q�L�g[K�jY\I4I�j;f��QՄ`��e�*P
�#�&����q��.�U��d���Q�J��R��ZC�Uh��U�����q6���5-j`$����Q]���w\�28e�6e��T���9~
Hq���A2BSW���L�����]��g�#5��o}I`ۺ<D�4����z�b�F}ѥ`X�+ I�Ƨ��A�l&��N��ZG8���$�`Z�de��E8z�����b0�,�F��J��_{�й&P�BK3M�
��$)��	c� �^�R��0J�*<k'ޢ�x被���$�aI� ugʌ�%�����$�����`�۸k=H�6�1����6�8���j%w(������Z%3Ӹ���6�iW�2�KJ�~r��b��qW�����ow�ͨ��EQ.}����Nj,��H��f�3���	)"X�4��MY�a^[��	A:�}���	ҷ��"�	sMpbt�d\Z����Q�Pv���x6f�X�j1���g4n�� ��C���H�
]Ź`