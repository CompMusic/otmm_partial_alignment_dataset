BZh91AY&SY��� ߀Py��g������`��  :Y4:ҕ�$�2��L�S�ѓԚhɣ�4�L��i�z�L�D��hd�@��L� �A�ɓ&F�L�LMDE#� OP4�   �`LM&L�LM2100	2d�)�͢�R��� �z ��xR��G�� x�l�+��Ip $�Ӹ>���o	��T��$��l�sj�F���m\��)JR��'�����������������ww_��I�݁z��=�U�j�SAE¥*B��#.E%v1D���%��� ��!�"�Nq2"���	�i����s;��~�+�nΈ��#=Љ��R�h�XD;��)��Ζ�	$[	]1%���R�4�ݾ�?V�g�5j$�U��Q/yJ*=�ХJ��l= �n	�(L�� d�3ll8�w~��7�m��*�7�����E9D�zD����r#�:j�'K�g2E@�w�!C��n�C�y��i�]��W  �57	��,_\]K_��<hU�������q�&Q9u�FNe"
u=�����ja6;I��B�Tj	1Hh؎)����qy��Dõ@t�Q�ۗb@�]N��S
[(F�`i������&�����M2c�b�D�~������W?V����:��ԉ47b�eLm�8�xv��üLvq��y��]>�yޅ���|R��T��T���"�;�i�q��uCį^�{�w��+b�2�mf����'i�W�Y��ՆML�p�KS%	~_��g˓̛ne�8w�Z3r�? չ��d�,=��Ϝ�	�56y,fY�a�n`���<�dGh`�Q"�Bq��!5��:ٕ���E�P.Db����g������
�uכQ[2�Hս��-}���z�~Mx���n�ͅ�P]8��7���0�h� ���l��-g�z�9�S#���tl@�����^{��SIf�0�$p����g��^<v�*}
�� ����7��X� ������=Ch��r$���}Ƶ1���A�@p���E� �.���d��	�|�������gt�sT�[J,zm��!�I+�۷���(�yP` М�f�n�^���L ��5I��b�*��j�ы͕t��Vʥ�͗b�-�fn�[!H��Km�k)v�v�l�4ެ"&��jɖ�2�IR��`�Ad�:Ι����.�dJ7�˜$����Q�ϋY��/a9Y��}�gk�����8[�=F����*���t+6w����T>Y�Rv��T ��ϕ2��㍑�t�4s �_� ���ڷ�ۑ,f�$� y��¯<��޷Z� ����#����"sO��G!��xA|�.��d=��~�l�=��Z	�t�5��]�W�J�%%�/�kPnji66�K�dA�A ��K�$��&��ҍ����Ӟj�  ��d��zb��ZdW�\%�ل8
AP{��b��vm�*�Ή�,8X@��h��'~Z�;l#���a�u�pĔ��&�&C�Z�6�,���-�o]n]��v4 1䭷��n�]�w�D�m? �zA���T&�� �sT�arX���@� F���w��q�i�r�d�-��@�z$E� }	�4q�a��"?��QU��q@ d0��P:p� �b���� ���ی>M�2�J9�f�_Na���<�4�C��B .���6u�@�P &|�Jx__N�8+�ѷU�ۚ5ԐI���tVg�q�&�Z���6���1H}v(��C�ڀ�K��S���i��x�;M� ǗM��W���  �Y�#n�%��x�D nMz,u�d^ ���� r e�g�a�p������o��#��r�@�f.�p�!?��