BZh91AY&SY<&z~ �_�Px���g������`ϱ`�^3�@��H@	���M�I����mF5�C��i���*@@   �2b`b0#L1&L0i�*��� i��    �2b`b0#L1&L0H��LL�<����F���� h���R�	
^��H "@I�M��;��d� x�	���>4@%x��Y�h�HYo_�������;���ٗ���WjꞫ.�32332s1ckZ�؈QI�}�U��11�*S�J�<�Q��o&]C0�!�$����8t��II���n��Nk%HȽ���VT�3�WK�� �m�"#6�fIJ�9�!�'5��]���Al�R��Kı�6E�Iz��5�A[�ٝ]���YM�K��๤
kB�V��gwty�� M6>5��u�n۴߿uN���|-��8/��j���7:'��j$Yć(��G*4�f�d�����$�Tܭ\t�9Z�=���DhGe08�Q�pK���'��zB�h��[�~XL�4m-��[�"%^��e�p+8��hT�"��P�� ���d@����r�Vh�!�![�1 Q��xo١`$jn>-�p�r��fz�@��W7�E��i�uSz������e�p��iIږYB8��c�x�۠6e��u�h1���K[併�#'H[�9{Ӌ�}r2T���*�adX��RrFp,���d �q��N<<3�=�ن�L�^��sT�YΗ�� �w��yZ ��`��`p����."8.�8�"!8]J}��`N�Hpヰ��0n4��q�Á�O �`��P�d�����-I�\�X%�r_�n��̊����q#�c�$` �.��n_L�2�&>�&��Q;h.��b��@���zC�%�×3��4T/Ūe's�q"V�z��Tr�֠[Xq-4ē;ʞOo��"F66��`��.�N�U�R�@���f�8� ��eT̷ �����&6  SؤT� E9�6�����R ��KYH��%�@��$���XZGqג54f���A�v�  b@$a��㯉y�^Qu�}6U��v�d������Òr��N�o)�Q��4'<8��Q��)�ю2��ޡ��]��L��=,��k� �B:�`6�a�@b���[y��x�{]F���J@�gV��d�r@���-�S*���Jr��Tb�ȃ�E�+޽+��������������*E�ثT�br��wL�XL��_[M�*4�c{��6��I�CC�cH�1I^����`��R(ʇoaĳR�/!�0���L�]B2]H�l7�*H\$��#?�9/��?��u�i�
`�J��{jF��0ڹB'�Qڨ�ǅo�JQ�U���a�PTWZ�GR��|]S,��z�jԔr�n��l���i��=�r�I!8ӎ	ڽ@�ˁe�W�H��o�1�	n![$�g �~�%(�%�����M䊪���pD$(b�B�Z�^�Y��[*'U��Q LD���mh� Z/ �$����Z�+�x֝(�x_��3� �%��t()pN.6kF	� �(�>H��_L�z�:)��&�9�ǃ=�3��A�{��]|��@���SmUT�����������1pq,��,��R.�CDFz�Ko��A�=C(����â�یK�
9�
:A�L��¶e�k�q�f��(7���w$S�	�g��