BZh91AY&SYrg� I_�Px���g������`��\ �bb�͵�&&	��M��F���0�M��hTd� �1  hɉ�	���0 �`�0�&���Q�z�&A=G��d�����2b`b0#L1&L0Ih�D�ySM3ҟ�zj=#F� 4 �a�<�`$&�؄*H�=eOrZERHw�#)�xՒ@�@�d�P�������f^�~|>*�����33#2����	Ԇ!�R�J;���z)�����
Ye��Ӝ,l��"$��ue�KT᱕�ֱ=�*��N�d�hq8���ߞMi9k��9N;��bb�0ݥզ82���K�󽩈 ���LP�R�o�Ż�\�\����n����aG`U`�Kʩ�j*c��ԒdɆ�o��_�nMaJ���a�݈I0x�0��A:`Q�%��%	�P��]� 2b\�P[㕽X��Ԉ3ŷY��A
���Xm-��\��6�ei$M�BR]���
��MƆ�Qs4q�d(BC�K�=6�Ռ���%cn�ECI�ai
�8!�A.쁆�Qݔw�)E�֭����M�TdM@\B�e�Cp�(�m#Z]R�E��ﴙ�C�bޖAH;&1��^��Bq7��rG�6�^���T[j04y��)E�·$��p�Q�`Q/�v�j��"/RrFD�~!�]�N�ڇ���L�ltw�Y�[7Ea���9L9؅ϗ/W,�7�q��L΅D����dl@G��}��t72�Gqb$Rɣ�cq��8��ޞ����ǅDQ^uUA (���>XQ:��f�2�RIU�׋v�)��a=�TFH+i��djB���X��.e�F�����j��CI�x&6�80���y�,Ss7�px����N�mkɲ��(��te���b湣�:�c.U���E
jI#Iõ�ul���Mz��ء`�Y�5��������-��ϙ�K�p�7��=��t�N��`�^#�$��J����uKjIi�P0yWJ,Y���֨D���� �r��"���IS�f���.��5#ʪ橥$�3�ljk��(c�N���-r>FZɬQT��*�&�B0�a���@A��5�j�u~:4�p�i��2\��V9�:�Lq*p4����f���V8U��C�!��K��F�K4��Vq�ɇ !��Y���܈�.��F��D�*g���&��T�n�۟���W�D�����[ԸJ/�e�$�Y� a�Sy���6�ա`��w�A�΄��)%�޸ ���m*C�#\��Bi%�d����E��� S�1T
$*��Y!�	As÷9�24oV��Y$�Բ��˘M�5K���\s��v3$�i�y4�X��K�(:�VV��麿9�:���q��A��ݴ�4�t��8-����8/I�9#��(I(���S���{�0��rCE�ɥ]ER��G�Ӊ�4C���ݫ��Tl��U��	-R�@v�,�%!=N�<��`�6s! �eth$I�Kq��R��Y�2F_Fˋ	�韐c0�
�A�$�i��1iX|x�
�43#�֣S�a�џ���X��Q�H���rE8P�rg�