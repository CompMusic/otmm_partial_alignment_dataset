BZh91AY&SY�\� @_�@y��g�0����`~X�{���y|���!^�y�I!4�
=�����hd��H1 �T�2�     aJ12�ɡ�L�0��0�0�JM)�����h    E$�j��2h�#� @M �!dS�)����z�4� �@,�"غ����_3�J,�Ĳ�6x� P&T`}���u�@��.��̒J.q&[kٰ�V#��^���c�i�,�˽�f^�31fkZֵ�ֵ���%�A~)��y?&�9KO�Zx��	���!S�\�D�Ql�*�z[�9�k$�S!�ٙ��A �!f&�Nh���G ��������ȍ�8���Y�fiV���,��B6����FHPe$�M��jf\"��� �L�Q ЦX�e����|V�z���`���a�άbN�1C��	Ϥ�����m�	�����Źs�ܢ/��1�a��6TD�LP D��6�UT)��gC<E3�kE0��m����S"2[�1�WVΔ�d@��ޮy�kGnCq�auZ���;0۴:L��0�#���+����!�y��9:��P����\�u��R�q=�{e�<�eB��x��1�<ow_u�2$r�lY�7bw������Ԥ�m�Dx���2��)v9����R����Z@	U7T,wf�1��gQ�l��� 2#<k`� 
*.@�"Dk(�[DP/.� v��|��9\Jt%�E8���B���M\66�y��4�;��8���lW%�[���axN�Ts"\�1G~�w\GZ�q�O�j
gN�Gak��_�~8C��c��57,S�0����� jˇ��=m���ã��l:X*%J{�SXV=QQ�x�[Ş����i(9aM
��0� ��i�=#�z�uU
C, -�J��
Bf�9V���ff[��Uv����hŝ0�d�	<�f)0�/�vv6y�T��LGn� �P��a#���3����)=	�2i856onk7f��N3��(�qR IJm�۝꡹�?���eɌڝ������L_֘��im�m��1@fYA�Z��[�����)k`R���E��`�Y���QTUj�Js������q�͏s��(������5lF����WQex]�?j��٪��9;e
�=j���t�3ii�O����-��afR�GJ{ԒBަ짏�Rv�28wA|��#>xHC`��
����)�F*
ؑ��ݛ�ʣy�3m���o7{\�����n��;x����~�f���������HWL}=Η����d���XfI ���x��<:M��f�H��
E"�Y8��6*�N�Eɭ5M�.�d7�p.5�4��A �Ƈ��W�T�U]dU�t%�Y��!�P�D°{�$/դ#��W!�9��w=��+�z���=�du��}Z�Sچk=��	փ[���:ZNY�����X-y:z�TaԪ�I!P���kT�����>����TZ�P5$���"�#�#�1 dՁbH_�j��ƃ)$t-�T� �[P]םl��L� ��P斒@M]XHy&8"!���`\+�N�EpO,µ�E.GKN%H�L`ˍ����=Ғ�Y2�5�$$����[v7�eb����3��~�|�H�h!Sq�e�,��I��Lb�ǹ/�8C*�Ue8j�ŕ��m5=F{IL@�@��0a\Gx�'[D7�5�{�����5c���q @u�x̒A��>�R��~��=��<3rm�z
g��c3$����pE'#=���� ��bO/4ׅN�I�^���YV��@JR(91�t�l>�V�*ׅ�f6�PI֎�Q/���)��l�