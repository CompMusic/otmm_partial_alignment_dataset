BZh91AY&SYAk�~ �߀Px��g������`	��W����)F��F}W��cǱkb|$�L�C*y��F�z�Ѡ�� ��F�L&��4�JyT4�44  �  ��PT4 =A�� FOA**y0�MD��=5    i� H� �4)��􆞠   4�iL����ƨ�*)2(P� �n�/�0��pMD<V��� KA�`f][����6m�O&�J�����s�b����ꪪ��ꪰ�v@�� �l �B��9����qbfL�6�3LĹ$�G������&@� "�fj��KJs�i2��2"?q�ߍ�Hۼ9﬊�	dd����Ӄ-��;�J�JD����a¶]��v�jH�������އ�%�TI���K����.'�I���g�#��
pBb�wr���ؐ� �ĲPM2�Z쀓M1�wǴ����F%�x���Po��E�;M��	9�҅A��PB4�j�#-����"V�r�>&x=c���ѥa 323C�bq���8�ٱ�8І��U������ ̸��u�9-(�oi)��2j�������靍)�/	�CQᡱ�rHK��	a��4H��И�Ũ�4<��J�����j�.��P,�����Z�E�ݩ�u�����=NG��L$��Q���s��Yz�+��DR�ؗ'��NZ��_�	����n	G1&�j�8Aˮ�ZD����h��ط'[	�ʙ/���H+
]���H$�f���P�e �ĊQ"g* \�d��,�r�����r'�.`�@�9���;C�w�T��T��X��:����Ix;��sZ7uba�g�o�lG�H�N��sk0�3�Ʀ&v9�	9��.\A0��MC<��L�P,�1�T!F�����PX�;(�H��G��Ê�iw�2@�x��i�5���S�Ad��E�X̷ �`���)6���(��ɶٌ��� c���2�IuX��#{�5à�h�X�\Aw�n-ƪF���d���uԔl��F��I�'���I���R��(�F�ƨֽ�,d�_D�o6q�|��t^�nj��{�"�����AT�;�}i����c�^C�U\m��.;P����t�kiX�eQ����w����0���udE�b5�Y$AAia%
�H�B��*��m��"�*��B��aūU�4�(�h���V�$�!�,�{!;[��=e1�]9��>p�=��j�[7<��JoJ�^�����V�<+���F�[k.��o�r;�P%ܦ�O=,�w���D9%�@��m�@	s��l8�,�4ʁ�NI�@��uk˵������ -5�TeN���UdA�A����MK]�A(�ul����~{֠�eA�񱪀�=ͤS����7�W��'cXU�Q؁[���P�j��k0�+EY��hsіe�9��!�F�~�3�@k�i�y"��Mf��"�(�=�f�v$Na v.�����4��׷� ��y9�A:�ۑ���5g�N7��(�T��ae�Io~��4�sI�+6`�ױ`Uv�ԯ+C I�ʨ�Ø��7�JR�e����ܼ��$���^|��L5�I�#TIZФ�eo` ��fBY4	a23m��R1���I�(� ���$\��HD�	c�"`%��)���ꊌ�2�O�r��Efλ�� �# ��f�����Y"���`<8R��krh���:��a����=��@�A�h���F���Z��[BPC��)����z���w*������g��38�u����P�~���?	�kt���Dc�P�A;Um %9V�qǄ�U�
��ˊ,7["��1���I��C�	�z�{6P��ŭ����O�H�Oj���\
�ޱ,�,䍨�����9�,˪1��f3�<�
�?�.�p� ���