BZh91AY&SY���� ^_�Py��g������P6����$DA$�&���G��y��4�B�M� ��� �     ��L�=@4      ����&L�20�&�db``$#SQ���e=�jzM4@��	Sgn�B�!�����I�w���1 � ����١%Q�:Yk�"Z�)�俗(
����)j��L��`b���egt4�wȌ*�X �Q2,���?��s�K6}G��si1�/b9�����/����i�� ��t��B���Iv�$�$l7�\�.J��ک9e~PǙCH��&��4 )��.���5-��]me��{R�5w�Te)Y�;+Z�GB ��2R2Kq�;�� �?r�]�4զ5�nikrd9�����JD2�d�A��e�$2� �tI$ʲ��5�asK"�"��F�(��B�|
�&j�!�I�3ZP���6<�L�,xT�U�:4�E�
��t)F�r�Tq�J�J�4�%��`>�SV�%���g�\60�x���6d�a��&5��oqjfN�^c)&4TZ��V�,��L��<���p�z#"؟ �BjX�Z�%u����b�����bm�t��JJ�+��92tj�_Kyg� 8��Al��1��(�|�0%'H�n��� B�4H��A8� �C�j�dQ�'G ��`��RqdV�(i`+Qh�p�0�V"*]���! V��w���SG��_Fk����+�����f�>J
7g;�� *T�6����$0����8.�и��L{w���Й�G�����}��-��54!���-W�MŎ�d3�b�� ���-BX|V)aՙ�I9���(���.p �/5м1���0< �R|z�{��]��R,���*R\~���wy0���i�7(Z�`�Vb�`A���Ac2N3���}��h�	���q�Q���^*}F��md3	�	��{ T��lX�����I��]dۑ�xF�F��\叮�zN�H�%h5�IDK��V6-ވZ�i�EKX�d��&��:o����W����P52BP5��m��L����!�����Ԭ/\�x�b4
�"n.��%&�/32gV������&�q�B�
��X�e��=�i�gu& ���ϟb��[tK���J||�w���F�iKX���w��~`����kωi�Bv�,4_�hbL��S���U~��*,m:	�4	8~��7lJ���O���.*�˔�� �[0����ݵ��q�M��p�_YER�r�n%6 {$��6�X _�n�����X��H�%d�(�@��l.Y�W6NZ����wG�c�I�4d��]��BC�/�