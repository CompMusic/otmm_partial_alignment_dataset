BZh91AY&SYF|_x �_�Px��g������`	?{q�{�>� �}��n�h�
�$�L�0�)�4�CO@ h�F��@QT2� �   ��PM1  4ɦC  MDB�M      @QM�z@4  �h�		1M���FSh�51 h h���!"@ � ��@@����qL$U���!#)�� ~0H���,����	9�K,����f��FR�;we)�y�����������rUUUW+�\mb��(_ԳJ�p⍞��`��u�F$�/R�!e�9��ά����JP��!UUT�E 2Q	�.JE��nn>�}�7��?�EJ����</��Y���:��C,/4.,��LVMb�Qxh���S� P\mE4*k�Q@+F{+�I���q�?9���n���C�$X} �Td	JRO,���� a�L�6FlN��Vbε�=J���1,Z�AM�"fIRX`�CRh�P��Id.e	�3��n"H��c�hG*>@g���Tk�!���,E��:�(��� �l� �D�t���JV1�Q���ui�X�)��z�1�%V/���PA�"��h�a*�r*]�r���EXV(8P=*x�%� �;(Y@� �0�+�sb���*�U
4�CD��_M�.�o��2V��0�c~��\a�����z�`3.��.쁑�b�h�ۖT�哀��B�|)4��/K�$B��{�ٜ�W
�����1���t�܉�B�pW�!때�9���K>�&m�q��=�-�U�6�\"�JUH�]�K����U��^��]s8�������+���Q�S���
.9z�qWb��ǆA��}��8R���D��TX�a9@d�} ���|r�Ql�{�)N�@��4����w
p�q��0-�ǜ��.�R�3��?�w��ȋ8�Y5[Mf����$j\�����NDC���bu"RꭩV(�������)5�k��m!�+QEJ�f5*�	u ��f��
��0�u���ߧW0;��w1|~SۻcI���/&�`A�|��3�f��U�jk��\#��(�%UPA$�g��CM|J)t�i	8��e}
U��c��+	�2)�/hj̈��QEJ*P��V�Ŷ%(�%@(�������Jf����Vi�Xb�U
�be��(ɦ������Θ�]�2!�:ӃK��f)e7:����t��
ee^�6pP;���2R������5��H�c��\J��5t���z��4Jg��m�1$��wb��4��F��d���r[�%b2� lH� z�s�V9�ʇjL���K_�ZBZ�/!�@'�s�%�x�-���.��?��=���[@ŐkA��3�Da(;��3����!��;H���u�	^uj�U��Ta)#�6Ӧ��a6ʰ�lH��V(��P�,���Q�A�
�Nw���2s��T.G�y�rႀA�Bq�$�<:�߸1x�S�7�Y������R8)PŔi	~��C�u=�JG�7�&@0IK�p$.8���MkUq�T'L	R����������$j��Z�$S�ƙ��Xͦ��K�Y�<�ZĒ�/`I0��������������~��oOf{<��@6�HKۊ�F�eKႊ�s�	w�t�i!,$��[c"�ԋ��K����cd
Q�rׄ���y!�����"ԬORb����RE*	��54ȉ$�L׷} �QrB^��Y�h4 �?�}|���s8kJ�A�i�|vl�%�u1�F�j�I[�$�,�3���(��jz:��Ӯ�EW*�9�͛)&�}����$��O^�~[�9���b��;�̐�d�s�~e�0]S8��<7WQ)��l	�BN)+ �Q(�uH��|LL_��$n�ҭh4�%�DmY�%��O0��� ���Kfk5�q�f��x%,o�]��BA�}�