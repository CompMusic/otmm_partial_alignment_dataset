BZh91AY&SY�:<� 8_�Py��g������`0���  g޳����v�HDheS��='�6Hh��4��HhjIOP��     0&&�	�&L�&	�����z���� �@   ��T�����hOM	��ښi�&��2 �HI�2���S1M�6S��=   ��m�ۨA(*%@C(�!�������  �@�`~Ҋ� ��p��B"$����{�������ǩ乿Sə��w�3���l^fe����^fe�%L��ٞ�p�j�AS��oL�XRʻ �h��؛w����2d���c� b�CBü�@T�UBx$��[#��ͯiﮨ8����}�֫&8�w;�z�R%���
��
,*�AbN�'�}��貈 �������6�F��.���qT:��W�)m�VV�(O=��0ę��m]��HN�J��K(Ik�f$&L0ٿǯE��v7{[Y�x�~9�LfPh,���Ȕ�x:ش<��/1��p^�p� R�!�"2��S����^�r���;�a�g;D�Q��kW;���p%zÏȺ
S�����Èo�P�R¬2� ��@脢�Ȣ�V-�v�f;��h��k�n�L��
\�D�գ��$kl�\�h,c=뗶q��Vͫ­�-/hW��W�da`Z�z3>v�E���@C���P�s���ޗoy�`�\G*�4��Ab[�郍L�yA�m��H��X�7���KnJ�¦S��zػ�NC���7'E�ę��1ܗ �yi�ڟG]v�h*/k,zl+�ph0�K��:�v��B�I̬�E�3��x�,_	�\|��s�z�����Hkv�fE�n�P95ɋ�ؑ�V��.�Vl�A��`�%�NՆX��%j� C]8p�^ɔ����(�~��j�)Q�pD^������=+ྥ�e����q�j{T֣��4����93}��D	�.�g*Ϊ�B[V�<�ٻU���u���8����+��
�\ge
T�E�]c�r�9s��Nh�d�Ǉܛ��pqE���kA+�޳d��<��:j"��Pd���n��H��-�X�	!/n�8W,��M%���cM1V*�R.(Je �"��Ō�(��U;�5�Wf�C	�f1l�E� a��*���CD8��N��v��V73N	�!��������U�R�-�kü��{g����}S�Ic�O3���U�n��#�������eJ&�:L'`�2 #R�6�<���8�GXztB�B�H*�n�8�����+��������U�dH#�&@��.�'�"���K�Յb���=W��3�P���t��\?�"�E�INbB��6l*툛@y�S]���u��4Ƞ�,""�EA`QՁqlΌ�\�u�fѿq2�I�:�2��d����3^�����a�KA�����AX�����Y��)�@�h:�6�#�g,(7�s�.���yFR��������H��aq�+��q�o�V-�B�h�!0��zf�󼎙������ӛ�L���(�%��0�ڎ�c$����2�<N�!�r��*7P�A�%uј$Np��hÄ�5� 	)��d38����a4L�SD���'��noR���K!���3
:��_v�Y@|����a���!����^�C.��F�/gB��t���%ϴr.���r%��6�͗h��������0����3��׻#����0o�N���![Q`��A\=/���fb]��v��Ѐ���
��4,�E
0���UF *��h��Q�3�5J�cP`T@���"��%̨��Y:�|@~L�V
[�����m�	��C�E���ܑN$8�? 