BZh91AY&SY�]�j �߀Px���g������`�1��2� �4ل%D$���14����!�1�h�����)�hHb   � sFLL LFi�#ɀF�"Rz=PѦ�@@� �ѓ �`A��2`�$��OS5M�&���� C@zOPi`/_%P���`�#=��_�dF�S�;�C�P$Q��T��w����|^?&�Nfc�&.�	�m�$��̜�\������#M�yVՇ�e��d����X��7�l��MZT�k@�d!#L�v��i�L=elk�eUЭ��"Q4��q�y���kuU��K�����w9?N;&�~�4��;�3���!�P�ׄ��� C��1(�8>|2B&a�<�-����8�~?&&���7PU��*K.�5QB�ukR�xT�%��U)Rwd��J��bn��i�~���͛Z�(egZ���	��	��`@ssݴS�N��P�xW:&��V�0@��B��R�Z
Đ=�YK�VMD�{B�.�m�w1��o�^E*��[qu��=T�P�V�����r.2�D���ơ�V*\t���u���J���$l+�U��K7Jʪ�ҷ�!��6�p�n��cTR�`8�;$�'��Z#�y9�9!���iLc
�"���Q���P���:��
J�N�&� 2!�_n��W�@�&
88�
���R�3�GR�Q940�jJ���nA(�v v�q�F����\5�jH�.�J�L���Y[�V�1�����<�1�uM��H�.�	a���M;�z�V� ��������ͥ�CS+k�]W�.8�iQoX�ﺁD��t#�6Ĩͤʃ�#*t�|��/`�Wn���n$�v�,��L���g���,7 UhƳi�Y�g趼��쐄���b��£����i�����7�J@�A�(�6!������^ET�ͩ�%E��*.9ܰ� �JDH�Q��R�UPZ��N�-<c�b��,a$3j^��߮S��ڹ�s��M��R����N�ns�}4)���5{��t���n��Bw&Bu���Lnn���2<!��v��HU��s�M`{h3w�۫����d�K�W�#���8�"�+!t�.|��Mު/��(�9�"�2�\o�)�;�G������՞߲
�
���d4�^���%`J����cN�`$�
@#�(b�`E�\�naܰ��c/\p��A�p�|��Ʊ�#�"4�v�ܘ�gTb`���H�Z0M�h�!�_��:V��0	CH���</�!�!6��q��|�y0_��z���ȫ
J�ٖ[^ŶZ��lB�r���ea���S���GG������}!����Q��A�#�y�&���R���v��=�Qw�T<��,7q
&�%J5}��o��.�i��nMك�3.��f`�3"�!l�E���I�?���/s{�WmF񙬬n���p9������N$*v��y���Dp��>#zy�ӭ�;�nLdeӗ��3�g6�M��m��r�����!�"��opxة��$G#96*ڼu�lb{�4�FQ��X�t��<�]���N�G��a<YD���m��S1F��8�G+� w�<(bS�2�>�������(��ܑN$;�pZ�