BZh91AY&SYj��� K߀Py���������`	�z�׽���@  <yL��Vځ$Dɢh&#�`�4bh4 z�h	�$�2�      "f� ��0 2d`  i$$�?%��  @4h`�1 �&	�!��L��Q&�hѢb)��I�?Rhz@��<���=L9�"��A/Gą ��|g�9<��PI `IP�s�
���/! �б�l�����q������^ezy��ZI$�I$�UURI$�ĝ$�Kuf��C�����5X�G�Ŏ��ߐ�S6�0���mq��hk��xئO �F���O7�qK��mm�v��&#�K�k4���ɗ3��Y�������;y�a��gi�jхmu@L9LlȽȊ�Pj���Ⱥ�ܩ��V꺦i�ֺ�ò�Hjw���( �T�	aUj8i��e�J�ʼe���lT��x@O}�C#��'m
"2P��۩�+n�뉻����a��<�os��X���ԙ���� �C����!������h�P@�V��Q"Lbbe��Q���[��m�H߁M�2 8����7�gi\�+��4`�	����Ցr�
�J��5^6v��˶x47�G �.��g�!x\�8�;4E����o�p4G6�xv"�I$�Ys��9�����	�&���
�d:��(uk"���M���כ�:׽o1�D��
O���@rj:����w�vná�y�!�hj0�F���3Yw@9���fCM��u�^�÷����40�L�<�y;��#z{��̻�9�뮺��y�c���@��LlMp��&E�z�9�NoR���&�"LO]gq�ʬ�I���`�r9��{��.�+~kW'oB���w��3P����qn\G69K_?Z֌h`8���W�=��t�V�z�Rw��I�)����D�tQlhu�
5a��ǁk V&	���wwr���P۝P3!ι�e�/���<�r����j��ɪ�ͤ��c!3Z�'YU�ͩ��+�ř�HО=
�m����Y[B�t8�uU\�xuwW����r�Z2a����^��+]�?n;<a�G-�r�~sB�
����)���J��;F�
��4�;���:���wyQEi]暹�x-�� Qy˟N4w��;�E��TPa$�=�|EO~6�w����n�$n��2���q�(.�ۡ��,̀Љ��������K�db���Q)h
.��`ȱ���
\j�fÈ/��[��]\vJl%DM�<ۆx6�>S���`ز2@3Lȭ��5���\��s�Μ�yE�^~�a��j#��y�_�E�=x�鬠�YVX�\ư&���~*�J��I���*���$�xw���?l[�1�?J�ܽȭɗ\�
�)*D����M۱�r��!(�?%ǡ3pL�R�] ��M9@ߕ��Wj�g�b ��|�]�C�
��P>��6m�j@���/tF4��|oҁ�u��m����ޞ��!���������&��"�$DX�Qb��`z}��l�o d���&lF/��:xKHZ�����
LLS�*[��vL\�&�/ʦA,��&��^ŝ����3�k����gI��N<�L82P�x��ߝ����ʤ7?\IPT�7䅊!�h�����i2��5��7.U�3d�+{�ҙ���@$�z!�54�o=���߳3w����c���� Ju����T�����	�\���_��Q	��W�j%¤�CHb(a�IM0*��I@�`�҈�vpC�{�BI�ٴ&��L��8�V�d�Z�t(WS��HL;�.�դ��*t��E���� �{��y��8��%���֗_xݡ�[��H�Q�5��%MJFCNn��^!h+u���Ȼ��糓Н��x8'l7QP�;��W"��X=���Z�o��aD0��f���I@��~}�୮F&�d���m
%4D��A4jۊ�[,e��	-eP��
�=���a������Wю��1�!�
�~"һ\�]tL�Z&��:l���A}�$?�N�3ʀ+ZS��rE8P�j���