BZh91AY&SY4/* A߀Px��g������`	�,{���   �ז܎�ڡH��M6�i�	�i�F����d	�Iz� �   ک�F��4    A)�"$��4�z�4   �12dф�14�&���2z&4iF�@ 2zO�i��=��`����HX+��Z������R�{��C��!�@-�Bn�,w
2ٔŹ/ӆ�g�ekl�k9�����32�1�9�3ff^g3ff^h���LE!���>�R��uPjH��.f<��\(��D�w�l[�!.��F�{�7��bK�a�6�BRH'��3��b)8/��<ݞ�#�P���6*�"O����D �%�"M�%ԢP�����%�VU�>h�LnϢ�G4�96�����7�^[�ٜ́��}��O���CƸ��U64�EM�� �G!8�E���k@&L3x�F�ŋ�gw������_%���R'�"@��z��=�1Tn,Y�K��|�y0 `���^G����P��}��o�<��"\���`J*�SpWS+g���v���ˊ�K_FM�/VO��t����l��Z�Gs�9�!6��#Η���{5��9U<s�Jݖ���v^E�!PÉEf\�*S�Ж��<3�f������t�fե����_uy����j�R�٣�Q��� �.@O�8k�}"Q�
��"��u0-V�igw�u���c�+�(Q�� ��1@r!��Ɂ7�[xr ���n��0�������Ig#�7S@`4. ��+ٽs={z��WG���l2h�$xƣ�ؖ�G,'θ~P=����^I�E>8�M�3S{Vޛ���r]����u�B�|牆Vc��j�h�8�I<��Z���G%(��g"S��R�CAeC��O|���~ՑHA�3Ĳ�Q�>�(sK�	B���*dkԅ+�?iO6�u�=�F@�py�]q���f�X�&�8�~x� !rJ��J% A�F��_�p�����.4��=5"� )��HNÇ}4�Y.��R�nJ�'u�'���jN6f��W�-��:9M�"�/+�̗���Ѕa�2�,3��Z�"�#�(�+�UT�&�/uq�����c��̠]��k�y�Aij�M���DR%D�`�h��`L44&R���ő�-(�$�Dnf%�L���61na�`��FI�B(�HIEs.֚Q��"h�a����⌻Z2!�\5��8��	�U�BMk���E,�ގ��O�=R����yijy��Xi�z0����4�+���2yK:�#�u��F�;k�]��݋��NK�^ H.ՎzA��w�i>?,�OZ4u��I*�ఫ�OOE��N���\��TXr[����|T�r�m�^ŵ ]���a�5��a�Q�� �x�<��.ۤ����G��+"%���*���J�����6�[�]����D����o
/�
QH҃CT��J���^UE���-U;4N6�T�1��ҍ����Щ/��ȴ��%��[#V��M�=�a��2)�~�S+V+�e^\V0�+F�|vIG��,|v�)b�.��\g_7�|j��N5I�SVÂ8�"�R,��|�K%�9��-l�<��v4t���:�5�����W�q^�k�7iӧ�S��k�k:۪Yò�Q����Y7ٚh�L��d��#b�s����UJY���Uz�._}D��t5��r�9�,�5�Ű0;L�$�U(�|DDmJ�*\���&�$�E��%KQ����9+�to��־���$`���@��[8�*؃������7`plp[�:/�w�%�4p���&~�1��̀��Ĵ[B~j�3�hsX�E�ə��`8A�	�������M���5����s�t�e,��	ڙ&�	��8�?�qQDng4���i��ƻ�� Jr$�쏓	�e������>R��׬s߶h�n���ņ���eѵ�V���UG'L͍3�O}[j�6��4n&�$�w�.�p� h"^T