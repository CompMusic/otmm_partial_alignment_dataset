BZh91AY&SY���� >_�@y���g�0����`~}�}>�<HF�x�m�i7wh�IёL�S�e3H�1=F��#@=CFA��&�� �  @  �H@�Ph     ����z� hѣM    4�� =M  4P h"!Sҟ�hM�Ҟ��țBda2`���E����� �K�|IE�X�����O(� P&T`}e��u��V�l����As]�r�������Y,����s2��������ffe�f]�4���PY���U�9-�4kU'p��b�Q�9��z��w&�7��Ny5&�"�A$IL��q�a��b^�R��������f�G�vH���M���3���j�x�R�`����m5ے�J%"N��OlEr��Ҁ��T�	ʧZW�ao��GB��Y�'u�C���\7�4��4�p$��ԋ����qܒM1�ӟ�r`ދ�e�C<ٛ z�`�L9b���
2B�]�*zuL�AH����)߅Px�χ�-��$�S�Ì㼨ע�N2ոs��A�G\�Rȴ�S���
h�����F��oH�3�A�C(�덐TijPԧ�! �L
O*�]B�%��J�۪(R���dXcTs;(��e��b[����b���5��Q�ax� A���C�G#mK����Z�B1@��SV�2[�(^�
HhxPHF�d'��s���:L`��),�/2$P6_Jֆ8̛�AX{	��4� f�s���h)8�/�
���9��J^C0���:�K�b`�i�{V�r-U
+��%**�C��e$+��2SW2Q�x�֒�m1.K&�*$�]l�����L�@�� �4Ri�q�U��Ȣ��b�HPZXb�zi3�pe�"�lJJA$�TAne��m�"�mUO#�����WR���D��	��iJ�my����oi-�gL��U`,R�J�����ߜ�f��g�):��XF,]�E��j��/������klL��m� k߯����V\����ąLB��[�n�$i���Yjlc	��6����#D(r̤���$i����(ZV��b��Mh�2�Ô#�Cd+\Q�fǱ�J˵� �[&� ��2��+d�~�Q��r��n_���z�wD������TV�D�����$ѝ�i�bxn�[Qdi�&nHá;�$��W���*������؍`%z;5�B�P(՜��)�A�}�`�_�bo�z���8q=�Gs�]�����/���r�A�t��\뿇!@�Lβ̱�7�3�Αu�nU�H\�&Ε�JM%�)��~�ƅj���
R�-Rе��FR�T3�@��Hh�q0�C�g1Q�K($�������@�&b6֘�Q�=k�+�.�����\���"�F�gCׯ����{&�1N�#Gdt���m�/ӗ$GK�z��fA������V��/IS��0+�q�k\��Fږc@$�W�	0֩y^7nBk���]���@��Ē��"�G�Q�b2���$/��j�����A��v.0U� �����b�&%u4 @n�B�S�HV;la$@��@��+Z�[��Xc��՝�8��P*Ȧ�5�gF|��Tq'&���XfHI�7�<��<gT�C+Ts��Q�n���� Gq'�a
��A����	>"9�1wx�UQ��i:xJ�����oZ��{�LB����C���eFwe���>��64�:���	wႪHVhz��|��yl�h�H�J��,��]]&���HY����P�x-�c$ٽ�J`�M�+{��t���FsV`�(:����a�7W��Xc_֩l��Q(Āb'�}�ܑN$4?��