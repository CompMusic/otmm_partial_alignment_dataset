BZh91AY&SY�q= 5߀Py��g������`_z�wn`  �F!M4I2bb�驑�z�4��4�Pi�h6I�4hED h      ���a2dɑ��4�# C �RL�jy OH=F�    9�14L�2da0M4����$D&��� ��O�=5���T/Ǭ@��.�͠J@{�!��0�Z�>t�I��HI��8�p�6���Av�����g�������ֵ�S0�*�����&"#'#/1�.��@�+�V���^)��ou.���TE�-PaT\1�xw��)p�J��P�xB0SY����n�{�H��#36v��;��4�°
Xaf>hJ[h��Zw��_���PHy�����n!2�]�/�y�^<��}�&#����Z�m��t�Z�HG9��̈́#��x�O�Z�q�V�z������2�v�R�Rv�إ^5��K[�`�c0,,��gs�l�2�#^�j��2�e�W�)��RT(\(���*�Uމ`������`��	#D�3%�C�3��G�vz�$T*2��h�(=	� D�w�w���
�E��D�J1x�-fmck�Y��.죲h�R"R�D�C�Ƭj�Z���n��׍f�샘D���(R��)
V�����f����@�*Ƙ⼯Ҕ���9�"�S�x؂@�KT���G"����A^*9�G����9f�J���E��?"dc^*��P�J���YQ�Q���)�����u=��3�8�/��ƪe]Ѥ���lj��b0ET��W�@��CX�Gq<��iٝL�f�k�,�.f-�yHC:�WT�ee=#��d�F;�I��*��en2�T)�I�M�C�n��؁iᚱ���u�̗b8dg��	ΰ�V=�36���c��9�wt뜎v���Ot�}c���u��v¨���k����i���R����Ļ����I�0Hg��OP�G����׍��N��mQW����	���&�x����/����Bb�qT�jJ�遚�z�1AE�",��n�,��N�HZ�D&C!C�tIf��)���L!Jee�̒��2f���υh�^�����pĄ�v���_�jh�$��?��zU0?펝���W׽D�+P�o='�G!��Д۱�L;swf+ц��WJ�Oz�Y�)0�J��R��7��֎a!P�np f@y�81*M-}E��:���C��;Ƅ!Y�[�f�K�^�\�����޾i��*t`�3 ��Y/*(�SL��'1}ׇ��T�y�z�k]V�D�qs9���B֞��U	h� ��,U�B�1TX�d8Y#�Ь
�ƑF��]�zK�D!xM �9��-��Z,<�5�.��6k��
�B��!��V�|<�ז�&S����@k�ˡKl�d�m�?�$k�~s��,z�uᘁB�pb��n���5�d�:�V�$&���}�k�E�Iz�W�Eٓ��n�!	DP�ؼ���r,�*,�t!'��6����H�7�O:�M�[N�$)S�:	��#Ƞ���$/l �+�Vy3�����U�N��"�Bd0��1��d�!>Q�5�PT!'0[�~0�7�.H=co#=���� G���j��b�!c��1�����B ��x�y^9xw���f�ݮo��fR;v�%���<��z�Û�~8�gZ'[�'J�eC��!X�<��^���ʔNns �3��A�ݹ4!@�F� �'Q��S�*
�Z�k	�i���S4���z���2�B�v�
C�l�m�����yF��#�R6����ܑN$8�OD 