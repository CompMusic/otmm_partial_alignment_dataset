BZh91AY&SYѵ3g �߀Py��g������`	����  ���i�A�T* ʦ&�d@�   � ���Dh4d   �����&L�20�&�db``j"�$�4�A��  � (����z�Sz!�����20�4F@D��i�"OQ�z=56���OS@ �z��i�a�T�N��J(B��oq)B$�H߼?�2F(� Y0)C�E�3iJ���#�0�B�Z�K(�� =p}_S�����T�O�ɬ�̬���l����[��̭"	{�	u
��0d&"Ip�N����K3*Aj[�p�ʆ��W�B��BU���e+t�R�"n�6&��g-�}a�H`0b��r��Ĥax���\6/�T����q%�I�(V�ԕ���[���K�uQL��υ��q�r����O˂����;9�/�QӰT>����1a�~�� TT��9�DH�HI�^��_��!�+g8i�k�/�ޛ9m�x:e�-b�e��!����v����x������^TA�JJA��mv�.��P����[Pβzr���R�b���*@�0P�Ҙ�gP6���ڃ�!e�kHA:Q�Rn��7��N�s7y�&�̆�s�ŭ_<UӔ��85h٘�E#](�B��4�_2��+f ��gP��R�8+(�^��]�*���4Q̔���J6�zL��j�R�ON�3��H���A��*OȖ���j- [iv�#�&"阙T�t���cj<	�&&N��:N��d��Owy��Z]n�$;b�a��x,'������0NC-汳*F�*�r4GB7#q�ޮoj$]H��.Yy��W��1���I��;��B�n�8�4X����.ؙ(��TҀ���Q�9,,�.� A�t{y�R�5۷B{vǮhS�A�BM��4������i�e�8}_H�hc�����ӧ�6o�sr�"���A@(Z�����uJ[L��'.mΙ��DY7QVD${x�ÆJ`$�0��Z�C�YY2��k��+~���8���B�U#�C)�؊
# ��g@�ȫ� �L��\�.j��Uj,�--�UH�ZV6U^j����.�]�$K��0�m
PH��51"��^hE.�<��� (�4Cev�<����4�^��G�K�Q��?���$Lv6?4$(�=Xӛ8}2�����8J�.%%jW��WP�D��q�Tr��@])��TB� 8�&�d0��	���C()�fbDN��d��''�+��z5.>i��������&}��3��7�z\M��%���/���us4a" �����C]@P�@.�'�1?<�k�`��
n�C�Χz�6#."��W,s��8�C��>�!�+졃,���׉�5�ǃ�������(�("(#�Q!�<B�tCn<����������.�?��rtX��I#"$�ዀ���B�Ԧ�����;��J�%��L�O��Q-�׫��ۨ����]n0� ����U������O���s��H���tBc��C0�'&sIXW��j4�G����i�>�?E�1�T�Hg�4������į���C?x��w}��h�{�O�z��"�;`��ZH�Z�5����̀�
�P�t4.x���]?]�(MF
�lhTn���q�l�t�
0�j�Y�Fb�%�@�L	B5�p�+�畁�B���faq6#�iծ�H���D�:
Az���df���;m:��t�9X.��L�bq�>M{ƃ��M�B�<� Tq>�y$��(nkIaRxu�^"k�����X�8L���|����ME�&�"B�@��h1E	�N�o�p!Y
輋��Y�6H�h�/�5C,X)�q��D��hj^�
/��z�����j�!��s��`3 �B�q�Qn8z�5��8�A���B�>�ǈ�vL����ߋ����f
of�_OJ>�ȯ�;��C�@��w��!�P|Ƣ�0�K�z���ܑN$4mL��