BZh91AY&SY�̛� D_�Px���g������`�,x�n  㹎#ZPH�h�<�JdzjP�� �i�T�04�� � �2b`b0#L1&L0JzD�P�=Q�h���b�4 9�&& &#4���d�#QИ�?J?%4ښzG� 4h؉�����֠��� %X��I~V" <�f�H��Q��#03$����ߐ��W�F0���~i�s���f�hw{����{�ʪzվ��'��_�w-���d(;3�K��TE�"���uB�ŶF;u�7P�H:r����|�1��IV�a�Ok���Щǲz��Y���s�q���Sh�+����8u�ff\���G2�Ir仲ccv�j�o������PKr�����3΅��c�ǎ���hߠS���.o��\����dиkaS��wlpB&L6h��c���&��.l�H(ig��3��6�7´e95�5F�A���@�AKA���>qt(�b�?bX[+u�f�5A�Ɣ��G ��9[�]\7�6�
� �A�6t^��%YNa%�`�e�w���HM,��u}I��.�2���n �"w�z*�bЊ	K��j��0����<�X&$@)q�#u�Z������Wu�!P�
Ԧ1�6�j��y�hL]�}���3�/��h��uPR����8�*��,Ժ#
TwPwYš+u�{��r%����`%�BĴT{0j�R݊�$�h􂷬�sG�!��ؾƠn[�B�����i���lM��i�ʑ�u��&{�p���v�N��.�"�D�e�)lj���#��e�ѥ��t7#sY�E`�*֛����mZOQ�W��H7����'�.m�.�8w�ݏ��~�P�t*����(�B|M�����70c����An�Hq�%[��T�b�UU8���K��o�o�s�t>�\Z����2��Z��;؀�Ȁ�����>�t�f�w�@\���=A⪨%QP���ׂ��GO����jQE7n�r����
�F�E){�!c��ah"o%;5��U��P�J)��fZLP���dTd���b@�.���Ɣ�%�Gh���{Z�f�u�i�hЅ,�U�p �$3���<����.4WW]��P:?�I|���և�����s�w�sTb�:0?m#���̸r�8�ӜP�/Jn��::�`e˪u�_���}"�i�� $B>�@��gφt�t8iP�1�D��?ƤG_O�A����޴F��}f�C6��4����$��	~��VD@�m�������%��i��0ng��	�.�ߍk���҆(Ut4l
��J�I���������r���&�.������.rM^]�O�d���4	�i�\�����Q�������Y�!w�B�G�y)gձ`���]��!�7xuY�_
W[�Do+�o�Q�J�[i5;�V�F�\�F2�unƶ���ZЅ�fa!0�U��a�~�����W�X�q-É$����	��9�$�&�8hb�����m!3S����U'�"$�(g�z��,�i�	
��o(%[HʄI30�-W�*��9J޵X����w�F���Ӵ�X��X/7��7"=�EP�xhh�����ه�ų��2�nA���l��nun�p!�3�qdQð�W$�DyQ,>�IoNظ���-�b�$�KH��b5��[Ut5>��lى�b�m�v�����mZ^��a�̓L����8��x�WQy|"?1d�m�,W-}v���5o��G�c�P���t"<l,��\(�D�(���!ƹ�'�nl�� ��<9�u���o��rE8P��̛�