BZh91AY&SY�m�� �߀Px��g������`
�,=�ڜ  P��Tͨ���W��i0�4L��1'��M4�Q���y@�@E)�4���4a4��d9�&L�0�&&��!�0# �P��&F��a4h�9�&L�0�&&��!�0# �I����&SdM3H������1�A'�X(�(�!�(:�E�V�"�b(F�:���~�"&}�B�d����l�����n7��Í3��R��ffF`�����̖������333.��UV]����$6����b��0l�U����+�ҫ4��ar��d���^�X8�b�B���<���5B�@
 J#[4��e-��VQS+!�mV	W�����.<Ǥܑ �ik��%mNůy�� i�5�l�b�u�]�S2�ց�������q��NE��;�K�A��aPS+���'�}5�ߪj��9oQrI��DM���:�N+G*�&���5Su�H	�M��*��qB@ɓލך���♝�򥦫��xaX[������9(��Y�U\���4L,u�j�-����l�mo,�ԡ��H�� .�6��]q��;���B؃�LͅU�2t3�]v���农
�0W%����9���h��@�`X�jFHuK`:S,�$��D�@���J�#U�%Q"���F/+�������1:q�Qa�n����e x0�*)�'���=�����d��0a]�5�{���Q�X������S�)E�*I	E4�M��K!eF�rB�Т��R1QHbUߋ�Q0Ǖ��W"��cc$�S-1��?RTVe�>Զ��F�w����*8�z={N���Y*^r"�%�ŵ�1\�4�Y�Q�j�@�$��+���W����7́B�8�!�ѣ`2ْ®sZ\�i��`�ȓl�����h+��,�X������e��nvq���F�[�|[OJNg��11�Aa��pH���u�B�49�(@�_�ݨ0��uF�����A�8��[�k��v��b�s�]���\+P��+�Qd������#k'QȒ�5�M�(����E�p� U5	��`�D9:�����,^|��<�G�����9m���r��n�k�~�.�dW)AO���5�g`;D�8b0`�D�r���ҫ��.˺is{l�:Y��nt�ik�6�%����C��7�j�)�냋3�"���j��X���n��El2��S�k;�5�P��%��3i �ub���cnK���pB�����IX���3����w���j"��U�Buux��Svyej���a 5��w�(EX�TTD��*)�T�1D�����A�S&!hZE"$UE��F^UE8�Ԇ!a��l�)eTPX,��ݷj(��Z�0i�eCt<��׬���40�Ϫ]���	3����{�������u�n�Q?hxJ�?���ZZ7��(���6����UZ5�yD��}U���9�9�zۿ���E8�	 �S��_Xh�i�<Y/�yEB���vQ:�%#���ƭY�y*BI��|-BA�ν�6��s�	�QC rh���h���[�{�!g��J�J�%��_��ˉ������?�ܽ)x�aY
R�
�� ����~���<VK9���1��pE"ł�*���(
��F)�H[�[G;R���ZҾJ& �ӳ���1�oE�(�!;ü�tU�	�*�Cե|@�lr�� eB��E�LZ�����ոw,A��+'|��]�[TF�@��5C��LW�Č���f�fKtN{��K�v�x=�K%�E�	��	 a��5~����!Ӫ�)ɗ{��;�4�.7�C��M���(:h^�M\a�:͍���ȦR��=Cn��g.���Ƀ���$m����@DW-�Ǚ�EU+	�9�Ĺ�s��G��R�yō��$���`���`�f�kBAǘ�,�0!�=���,CŜez�Q��h.��7�4����q7�AN 8p�f�M�P�"��ts�Ɂ���I�a��;��b�vvMš��:��w;&��n������J��J�5	ڻ*BA"���3-r��!c9�P@,��u���th42%qj�Sk%2oYM��-�`�w��\h��Q�jBA��-�lb�H5AĐ@ۭ�~�dN�[}��"ꦂT�,6�6qMEܑN$*�y��