BZh91AY&SY��HD k߀Px��g������`,=�b� w
�Y@D�4d4LS�MMCƦ��򌞐��I�4�Ԓ  � 4d� 9�&L�0�&&��!�0# ���H�z���    i��&�&	��0`��"Rd�1C'���h @i��PW{�"%A�D2
+?>�T+I�Q� }zF������@S03 .�&Ybom���D���FYJRʖ��n�����2r�����_\\�'�ρ��oغ9��	���~�a�����-dC�jV���5B��i<0R�/!`D�)d���2y�bH������$H� ���uJG��'q��l$p�ۢ�Lv���|�u�HD���$"��z�S�8ҪO��vb���ᡳ��,�ش΍$*V��ʴD�p.4��2a���[�>�W�M�羱]���
����R��F��Wn��㫖:�F
�	+
.�)��d��n������4���!��bɠ�ô�4����c���g����y���.4[ЮWdf�q��:(	t3�G�#�ׄu�.!1	Lo3FSN]Y��d5f�m�Ʈ!�BfK72�n?/_@�ű�pG<Y&R&L��-+�IԶ���!����:�"Y���J�*C776�0���I]#� �^���)4�(�6@���U��b�bW�4E�D&�Q46�̶��;���N9��&lS�@�=Up.�܏T �l26�����[��(��:�D�[��/782]�&" �1�F��G��:�hP����L�q��0T0�<��xT7u!�Q �5�i(�$���W
�)\^�e���a�� �������W8��e�6&Ag*j��ƕX�i��L��e�E�ΪGDfw�j�7�D@���>~�ouL����]{
���Rn�ܴ݆8�к�2k�� �
pN%C�xyVC��
�A�Y��J3�)I��gft��lcco���`�J�~x{����LNJ��	J}i�;���0l3R��I@��?���`�+zX�"���m������-��1�j�L*�CnC,
b$�4�����U-3ı4{gZp�AFC�������2T[W��z�ǔ>7G��Aj/i�S�6�ܾ:O�ziTVOT	�>�O|�Y�-�PA����K�[�	q2n���d�a��K��G,�!����g	,�M������M�fK�+B��ԇ�����w��G7��udB7��#�� :����gc���n0�ڎu�΅*�+�9��z��ߧT/�4��.�6=�o��n�y� H�  �`@�H��h�N��es�_!Z�s\z���X�rʍ�p�J�搿_ڜw�]�i	�9�Hp=�T1Tx�Kh�z������0�)�(j:�-MҎ����S��~RU͆��<IŞk5�?n��LU�Ť�E�l��ױo)�~T��!X�0	0ٕ����8UU]��W�3��f����$.���F��i�Puг�w2��6��4�4)���@=Jj#
��F��.+X�'(yq�(E��$�I���b/Qh����!m�L��C�bYQ�a��n �|�$-���~�n.HI�?��Hx�^�,�z���u�vk�/��r jM��mNT� ��ͩ�Q�Tmc��/��#~g7�tU��2i�cn���A�mzm6w�AnT�c��;��`·J���'΢��bm�I
r��hV�1����@2����$I�B��/��������n� ��nD!ԙ	!n�$t*� ��F����6�c2<�
z�Fo�c��PB�ap�?�.�p�!O���