BZh91AY&SY�E�( �_�Px���������`_}��W�w{� �|�}�R�mW��H�I�&ɦ�OSSG�dh4��F�4�@       5=M�҃Ԛ@     �MM$M�@�    �&L��h�� � 44�D��m ���4�C�ɵ  �4�]0Bx� �I��������K��46��4���"�Ei��,�Gd	N�e�&����}Z�a<���D�)JR��ffff]����ffW ��r����Yz�Hj��bo�6/G�bh�wNX��͚��v�kED£`�V1L
�0,a0�.>�
^��'+��F�+_���dZ|
���t[K\�j��0�Hb%T����Y%�=Б����$�	R�U��4��㊰�t�(����kW�����98�S�gq�HqH$�q'��t� �ƛ�xv��M����Z��*B����<��sE2��W�%�ɘ�q]H��C��ٓ26�΋nu��F���0{�	�Le�a�3=�fh/��rV*�!Q�\;��2�,���N�c��Z�����_��s�CZE,��j�e	��,��-�	B�ul5 [�Lp��%�k�2�F�rX(�ˍU�:������gY����A��|[��@��(I��ETT39n8W��#J�qv�RBR�YG!<�tϪ�\?,Yn�*_qc���`f��Z�(�� ��T<k� VS'QYG��\=�z����u|5�Dc�s���v�TB?z>&K~�&KK��0r`�fH^���S��]SV&]�2�d�	�́M�x@�ۥő >��.#90����6��Yv}J����?(A8p��م���\I�ǡ"�0yu�*��'���-�{^H�R
x;t$�|.�< �
ɏ��(�z���C=�Vn����uQZ"���~(����&l���1�@�� BI2!s6����w�������U$��V��
�ʟ�RX � Z�PC+u"@Z�AD�5�� H��H�6	!Z()A4!hK���D`�Q%B�T�Ĭ�&	dVU#�D�\�u�7ƭ	j>���f�bL�za���Z~��/�E=
e�q����x��hh��PS5�+^��?�(Y3�w����!���ŃWqa)K��~ ���$�5�ұ~�w0��ؗ@�9� �$~���2��ڕE����&d@���$�v+�bӿ W�v-�Z���ɤ�~ tc�F=����%����u��f�#�iE16�N�gSw��)m���J�� �S�I��6�F�߳�����lX0l@؛AB6�@�����,i"g��ӝ\Q�d�Vr�(�:��\4�I#8�fvI<=ek&֙X��>J� V�5�f�t$Na tI#�Bo*�Ե%����� )���NL[j6G�����9�_Y�",�I"˟�����\�52����ʞ�����B�$��[ Lz;u��Ԗ5e��k�����������d�:���2.�`I+\�ʌB�?F�n����v ��1��dtXH��KA� �X�稐�����vWb)I m���Vޮ���bȱ����'����"�C�A���X�)$o���n�@!C���� �8ιPxM�m�C��p^r�)��MI� nL0���^�Fб$��=�Ž��9��� ^:-��ۚLa��h&gޮ!�&bTc�
�
�q2�����
�<�DD1��'�,����� ���~R�s��*�H��R	�EtE�(���<�ؘ�'���3�sA�$�����ʔ Zd� � 8�{h��*�3%���7?��Q�
Q�����"�(H["� 