BZh91AY&SY98�# d_�Py����������`	�z�wG� 4`1ϭ͹,���В &�?@��ژ�)����2��)P�`     dɓ��&	�F�!�I�S)��hz�1� 42��55?U?(mSz���TmI����Mhd E���MS�dji�z&�44h4����T�q%�~;$(��^B��̤Y$�FQ��<��@��^�,��
�B�x�u���Weu���mUe�wv�7�w�Wd���f]��Ue���З����m�D.�?���8���lv�A_�$�2�q%�ߵ�%aó�=�I���oe�I#	�m��kX���T�~��ΐ$��bY����Q�.x��d��M U+����J9���P̖c�#�1��=��r���Zf�9�}��ǅ��T�%�ٙ�M�F3
,�O",:I(FU�8�y���ɢ�$�&C����#/�|�@�7i���j۶0�+jAn�0�)��ט�L�i"���H��Q�L[��մ�Wj��Ԣ�Y֡�vn�A�iV+6���F�HdDD` ^ha4���3Љނ�$-Su�Jg�t�x�$�II����2���IP	�AEU�W~���w}�YݰU $$�P('╕�r��c�L1��Cd;��t�Z�Vr��w�a���\����]�9:W��;����6v�X�b`�-�	Ob)�+"Y�+��P匽� ���B�rt�t��C�1Ҡ�5�UԊ�R���q�g��3mY6�Ll�( �����+�&��X8�e�V!��E��{�w�;`���[%֨M�b�;@�@8�ZW�Ő������B.�a� F
G���΂�L^	`1| �GQ�Zy
h������R�9WJ�V@��+[��1�,�TCq��;����7|�RE��R
W��je��; �.��*D����*�*�M��ɯ*GW;� �o.4]��)ߠ�q��L��V���4�`U�t&҅;�4T+C�JG�~��M�$�l�j�v7��)��P|q�Բ���?��Ls���uŁQ���@Ņau����vewyD ��:Q[T��WX�]��,��Uױ��obDp*�b�p�ʔ�I��v�k��ǵ���+�FI%)�]P�Hoߔ�}X�h�$��z�Y��
�F5�kKQDkZ�R�e�Fj�Bi�Ӝ�*eL)�2*�6��d�,�ʄV:�&f@D(��(㋇-��MEQuhim`̎���q�N޲M<�i��,st!3f*ȳ����J��c܈��;��B��џ�p��������Z��]I�iD��_J����n���괙�>�T x�>δ\WA�:��"x[��\�1v�� Hr�w���f4���t�DK�����N�ø~��L
��/�����g�o�"�oae���! %�v�\R"�%0�:=1�U��m;Pa�B��5;�$��E.h;T���K�z��$����
E��(�DQ�PDI����s�i�Y)4�$+i�e.a

����(��=�&9�U�,��>��c2��_���0X*���I5�x�Ǚ�J�7u�*��
�YP�<삑Ĝg�;��hJȩ�����H���,-#�:G�q��(pr$����ς:�|R����r�%��d�L6�O���w�ҥjv2�\�~��Q�}u*��o
�.�!07��֩��*(��p��kwl3�7��H�FiUo�n�0����$�a�������	����Kh��HK2'A7�stA7M|��y��{��$L�ّ1c�hU�~�Z=X�\ @t��}�w�C�5���L�H�p���/!Q�����*�≒A S$���fk���+�ǌ-�gB�iKҸ�1=�ĄHA�k�ܰ�qM�m���y2��'1"Y)��/��R41.ċ���n�p�cRa �����T�	%�I�}�� ��ׄа��mw	�W��' ��d#`�n����؂[�.�V�5g�7�@����d�Ad� �7sQ[ř,덿�w$S�	���0