BZh91AY&SY���� ?߀Px��g������`	�{qٺ   @gR��Z��BI	�@��SM���䟥3P�i�<�i��Q�� �  2��12dф�14�&���H�&�12=2`#&LsLL�4a0LM0	�C`FH#PƉ���45�L��\d�b�v�2�.!T�Q%X��</��d$,$�
�x�0�}K�� D\8�-o8﷏Mr։gEUNs������3kw7e�n���������ww����v8���,���/���𿧢�E"d<���!ש13�[�aI0�����.���3X(@(~y~�e���x�Yk�6�U(�B��rB+t�;ڈlo�WEB�������+ߵu�SR�v��_�V{�|7I�N��}zJJ�u�vF'��`/k��Q��c���{ݹ��/oj��lu/�|5�{��&;��=���&!<')��D$�:Kg�>��D#i9�Jws�/��Uv���S��<����<9b;w�e
!�ǔ�"F��P�*�nw�z")j"��pG�X���ǎ+��9�U-]Pџ�6c�Wg��B1u<k��=D�eP�L��#��F�?7��OV,^��a��si�:<o�[E&YD��i,:j�, �Ҝ�D&T��B�}0@�% [� iW�gk-���}O>��;US~��#���C��5����Ռ~�4�A��"��W�D0�uV��7�KQa�q�!��o\����&��(�]E�{ۓ?W"�s�#��By{�K��E��%�˓�sf`Y��10��/�r��w�>9�mt�"Ldl)Q}���N-�o;�d�!���G��c�m�dO(QC�Fq�B�8��@�u�Pnޞ@"F�P��V�
~\�FN��(I�R#�	�z?d@��4�_|�rqG���#`h���t�m�k\q�e$��{J%ovE
-Q!�*~�iUU�\9��vE�wsj^�0r��M[�΋�T���
� 9������#`���dWe�d졝���N����:��7����^����C�=�n�@�����
�}�ONV/HI:�u �S�e�U�T�fgUA���{O|��nI���O2<����G�Y/�y�kɋ��2�D�Ӂ&�M�4g-�2��g�*'���Z"�����U��xX�D̗��Z2���P=�pE�D��RBVh����ju�y!W�X0����xi���SK��&�� j���J��eT_�B�X�ܶ��t[4�#���)��
�U�b�K�+�#p��II"�%- 𻐶Ap��vM]vY��Ub����<6{9�2����/'5A@���Uɚ��wkG�(�W�z�|_�E�:H}�.�ODn7������46cQ#���Lu��N9�M�أw栣0H<�n��x���?����Ҋ�tg�P��l=�����}	��uՂA�m�f��Cna�~V��^�'cY�!k��j�d�����T���ק����I~3���������V���Q�N��4y9�0�{�K�F`b��dd��bȚ �(


w������o����=[�5�(�,"3'���ۣ#f�ɷ+�t�ApL5�@�#0(~m%:�6mS�Y���I }�\��s���M����aK����@f���PQ��U��&/�Z��IO�Zk�B@�^Z���n���?t��1����Rh�(�
��Bp�9�A��$c0H>��Τ�	u��dF���*��E�
�Jg(�8�%����!I z�bM��\Ӻl�v�mvV������P�`.5؇>��90 �+��s���9�z`��/�fi������(n(g!���je1�!�A	�g^^����"ïq_>����#�۾fK"� �����7e��"�#�Y/���Q/�Bf]�v���$������˅���l]Z�R�<**`HA�p�ؓ���t�ݞ��h��/	�b��0,+Ç��1���E	t�&pD��Wl�!��7�rώ��r��EZ��H�
?��@