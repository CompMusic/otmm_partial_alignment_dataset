BZh91AY&SY�6{ �߀Px��g������`�{q�&  ���&�*D��z�I����?$�@F�h4�*P      �bdɣ	�bi�L#0	OH���24C�6���FA��F�49�&L�0�&&��!�0# �A4�4<@joRh=@�hF�,��OO�Q,��Cr�Pw��>�ĥP(=`U5�[�Հ p .�!S�0�&����y�;�c�R������jS3'2�!�fffff]ػ�����} �S�[oԻ����ӥYB���2%D��a婥!f��#V�C���C�VVv��fe��q�.g�rk��T��?�[Y��_9Ι���\�ƘN��w'Fs�1��hd��E���c.!xAg4�8�EVWi�7���Lge{���ڙ�o���e6�K8�Rn2r��5J�m9��~/g���a'9��|�����;���ny&_?:����!��.��]���Vt�l�r���fHmJk�PU5����;�H1�Rm׻�9v�r���\\���{R1P<DX�@Z��!�� �k���ʌPJuQ�p6]\I|D�5�bjJEƸ�rpf��
�Q���&%�؉��ˍp�/�p�Qr5D��.�
�����ȫ{
�
$ÓZn�3X������H�g�!1l�+�P��N��^q, *r������? 4a���e�D�S!���
��`�����Nun���9	F\�X*;�߭ +��q�Wvy�a�$} BT(��u�3���I|�\H{q<\M�KV���,>F�>"u�	�%&9{W���I��#�ɱ�B��<2P�.Hv�U�bF!�6�t� �����)ho��bs�[�1�.�K/d��_1�͏ �28F�-�"��=3�;b�n��D�����<d�vy�`� Dy�����8�σ����5�T&������sYxl�B�^����X�[�Ӛ�I�5EF�]����v��g
#sg9I��Yͭ������UA��`�Ξ�}Di����j>��f�M۩޸}(��Z�}�8`�9%o$�8�n�E�wN0f&3P#$�D �j���ɂ�d �0F1�J��i]8^��d��ƗME.EVBZ {��G�{%�.@�=��:���Vʏl$�x?���W;����B����*?2����N��K�x�8�iEV����'���u�:i~�O�I~�ܨ�U�C�Bu����Ɨ2_����b�G_E	=e �^'ź��ٵ���@��a�p	l�}�9���]� �x���ⵧ��B:9��d��CwU��fٖ$�V��u��n0�Ϋm�!Bc�UtS�	j;0ŉ��	0]��{����ju��EW[\�)T�T�`j�%"������s���t̥��ڦMSog����,}�H�ҿA�˫�n6)����uL6
� Wڡ�.��c�-��0���$ �[r6��S��!�`F�8K)hz�
��$k���t�:q:���`n{V�2��,�J���a�&�j�b봆�uj����*�q�/d�JH	xh�@���<���B��� ��ˉU9^��9IP�*k���:�^�9�а�xz��Q�� �KI��xQ�깷oXgz.��e�̸G3���g� ��(=��^���ܹwP=x�ާ�˝pA�`����h7 ������<O9�t	Sp�
���	p	 �O�[,�H,3W"l��I�4L�7-GW�H-���_�׃�c�g1�\�g:�F)�ۨR,��8�Z�-��Ș@7�a:J�tJ0	9(b�B�M8x�So|�� ��=N���;� ��%��T�+��h��F�d�JUC��zr!ҟ5E�U�;����"�(H\=�