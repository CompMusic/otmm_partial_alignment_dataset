BZh91AY&SYN��� �_�Py��g������`�z�k��$  ��6�3��D$�##BS��2zS4F���MS�Pi��hT��      �	���dɓ#	�i�F& �&����MA��d� =���&L�20�&�db``B�h����� � ��	+���I�HH���	( o��T�&*��	H~���� �w��� ��Y�g�u��}�9�۱>|ֶK�c��ffffff��ffffffff>���Ç��LAo@ ���Ap�#�����͡&��[�֢�J�s��J�Ц�0f̘���Ԃ��¸^��kL���c]=GUk
�h41,o�<*�d�S*�2�CC�-�S�bɄ0��e�1�3��s �mvP�^�m<�8�TOm����}��F�JfOL
��V�SV
Ё�l�T����U��>Z@,0��z�x2��'���=��HU{!�l�wt�'"!��P�R���+�kC���p7=�lVO´sL^��//����j<�D��	Z�m��>�� nM��'%�h���;0sn�"�4�y��M`�L.�������abB�8��=�|�!L7eqؾ����y��.�#�uķ{���:}���S34}1I�M��'�4[�X`ā�<�Z\$$��1"g�i}�P�?Z.�"��Q�B����֢��޹�y$;�,Ibw����l�E#�q�nh8�	1����E��`.��y�k]�����ȹ
[R�@M�:�j1�&�Ͳ���3iAw�N�jP�	��1�x`j�x��Z��6�lk���:c��L08�!���hUf�J<�!ρ��6�`��9*��!"e�����d�I�N��Ó]�c=�;�؂�I�6 V��.4�_s�{��̽�ZV�5#�]S	71sX�Z��3�O\~Ɔ�}n��1�<.��t��h(��/~�d��ș���P��Ⱦ@��KX�YY�jx1J�3�9GV�اb���؍;!2��u��C+ � Y�S�V`CZ+������6=y�u����E�UT4'���>r��o����y�$n��e��E�UM3҅2ƕڪ���e�-]��b�QDb�j�*ҋE�
l�U��l�K"!5�k�a����(C.���V�
Cd=,֙��!���qgd��d�M�«�k��.1W���:�A󟺛��cʜ�"�L�*o{�>X�Wr��f��GWK�a֚]����K��ʀ��G�Q�hˀr��_*޾��8j�!	�$����eu�c[,�~�4��r���k>��=����t�ת_6���:&�7��x�{��M��A�u���f��\�\ȭ-r� J󻑭��&��n��N��`�1$�*�`)RAH�,L���skd�1��g��r�w�\XB�� ,�D���]�;&�X< ���A�Ĩ�SSL$`�_q�?���\�A����K�Y�	����-��WC�mٹ�n�%U'�{I�H۽��9�Q�V����B��ϞW�yS·`h],��5ӯ�HG}����m}��kr�L�a
�I��7>�!6l9J�ŭɫ���K�qT�d^��t��]W�s!��#��@r40 &l��^>9����P�-hj�Y'�S�H2m.i8��1��6��m;��@�0�ο��p��HѴ����tVP�=���~/�$C��!��)E���9������gv�M;�9��gH��2�ޛ@]�e@-'��U������sn�÷e�f�Lp�84Bfq���:ަ��٧�>qE�5ҝՔ�MCf���͉�ÖN8��U0j���P 8��R��p�s ���i
VVh�R�o�E�@���gH_F����Bz�&�%��$	A�S�<���6)Պڣ���F9_�Y�h]�rE8P�N���