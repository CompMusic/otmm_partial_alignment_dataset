BZh91AY&SYm�95 �߀Px���g������`�z�k���.T���	$������z�ҙ�=O4y �S2�M $��@  @ �101��&%="B��H4�M4d���1�� � sFLL LFi�#ɀF	"m�MlSG� ���M@a4$��w�����! �  ~��֘���
�����?� �x�;0l@�����}Yp!����w:vֵ�b���n��.����ff^fe���6[]B��K4/���ˢ��bI���D�魨�Q]�V��^�슡h ��ˊC�˶����CniՖ%bC���_�m��|/���	ff��Յ3�1�FeVf�Ͷd��aw.�w.[yq���䶭Fg^�Ԕ-ͧ�@�^��	
�}<p��Ż��W��t�ۼ�.�ZC
�-�Esr'u��k��#Εx	2d�7��F��R{+��WEVS�;>7{q&m$��Y�,f�B9�2j�B�*��ц�T���h�3k��|�c�@��� ��q��A�c�j *Ru�<}("�L$�Ɛ�0��2j�A��q� � �ˇ%0R(��:vQ`P9A�Q���!�
*&��$`��U��5���<x" ���A�T,F��h�oXXe�P�@�d�}�Y`
+�ns�H@��� �[��B,�
`�Ys� γȜ���x2e��6�Y��[�!dc"�)�"6Ki[��h���`@gRN�*v��nrjЈ�E���p�dbĺQL3��	u��g�a�����IB;�	�|�Z�niq6�zbB:�^<��8��"��^�������0A1�$ْc�I.4j��j���T�c��ZP+c
�Ǎ������*��G�x2��Qn��0��jE���p�ذ�{��&��[�� D��i�p]Ox&��5�����k�E�+�7�q�E��3���Hy�n�N�x�SQ�G�T�YC�����i���%��ٻ ��%�m/\|
�fŌI�Z�l0�t��6�66�m��4	8'OO�^%�MG���*�hu:�W��!;;&5�.6�a$��p�5NJ��P�%��� ��E�a��J��Ri�$��R�E�U�엦
���c(Ԇ�Ӎ�ۥV���!��w��i�B5���m m.j��T�����|���x��~ӏ��������ڜ���/��ֿ,8T���#�����r�L����<��T�l�����.���%**d�6��@�dwm��32�|��6/S��� %nU�19�0�}�o^��O�
�q����TEȃ�A�,���ہD�J|�_f��)|-�9�ZZ�Z����FV;���RG������Hb�u%�@�P�B�pH�Tj�Xx( 4�,�7Lɟ$���=|ME�J`%�lhD4
%�֫њkb��WZ�X=��l��Ao��u
��/���Zy��g������ �%>���Mdg����ʠ6�ʘ��@T4&H�+�ۜiˌ�d�MF}!�(���_������:���?MsM7��j��EL�ID���/Xu��DCF�(�Gp`^�j�������Ƅmm���3�K&��@Mq�BB0��Hr$8" h��%1�e56^�fO:
�i�L��(L�W]��B�TYm"��M�BI��ѯ p�n�猩Y�h*s����p����<�p�^�S
r�� �0¹�E�%x<�wj#Ղj���1��$Q�ۚL�Ȁp��x�8B��CO�Y�xT[q��]�+��(x�p	P�|AK"x�ppj,z�q}24�SPH��@%Jy�t������d	sM�<�Z����[�[޶d`�.��h����<�G�ҩf]Q�{��dO�4�h(�b��rE8P�m�95