BZh91AY&SY�b�� ߀Py��g������`?3�^�yH��ﾯ��!I0�D&�`��M����CMH �P jjIM ��     4Ѣi4�h�      )�"�A���@�   T���oRd��#M�i�� D�Ѣ)��~�xL�I=M�b��M� ���t%�D�h<���~���!ވ��nU������U"S2b���;�N��������$�I$�I$�I�X�LI�8������Í��� �nq[��D�.lnmV�Մ(����XiE�Z�q"�/�b-���~���?�����lLm��٥hp�C��+�#.e�8����
���w	�+3�C����`��H�k��	J�E�~�mP��W%Q:��Z�34F�����Kgm3Dpn�؝��iΈ����n-}���d7߃��U��b�ᗁ1J��L:�.��P��B��'l9�<���&�
��-����i��S<�e���á[�&>[�G~CH���G�U!S�ht$=ӇA�w�a�ä�'��vD�V��ɋ�q�_:��a�_J���:��X^��x_ �Շ��qF��[�U �`�p$��z��&�ȑo�l@�B�� ���v�X�[��"ʩ�[�(�Ki��K��W�-K�X���"����Z� �/�̰57O0J���Z`+6�^d)�F����z��i�8��bu6���.�̓1YH�nP��*��N��R��9}F�]M��������kX��Zg��
��FՍ�Ϙ���*.��kQ6�܅E
"��pb��u���U��
��K+�r�����R�h'�q*���*e�
�`$�i��>R[����C�D���q��[�u��-Y��k`��6j^�	f�g@/��P�}�Uf�q�;��\���.w�K�'F�B�R��f�}��Q��J+�8+-�8�j�E\Ʒ��}��:*"��PJ��&�g��h�+��k	TT��q���k�LY�rȬ�(H&�w -D��-#T�@����T��H��GG-`bA&[US0��T��VN\9r��%��U�C��D�ge�h�ַ�mJP
P׸��]�Y�uw�z�n�{@b�<Q��9���`��\��X�0p2�"���j���-�v'�B�)��8���y�/�����" r�������<l��i<��!
�Y��+*����eѨ5nN�R��Z���(�/a�\K�}۵����lϯ�*�o/j�����T�`��W��D�" ^������R�((*"��
�*-d�q���C&Kє3�Z&!7��L��"�!��.���/c��<�	�j�
�p�>���|���5����s��h��z��?E��6��C�;��yȁǕ#m/Ȉ���Rr�WTn�e%��"�S����i�lM�q�l�I8)�l�$��#��{�'�"�$,�P��v���R�$uX��H֭S{FAW����Ŏ��,M�J*�
>�l�[�pʼP�Z�N��˖Df0�����&�Gv���B[����ҕɻFT��(��ip�a�	�(�G��;��:E��(���}IԈ��8����Yy�8:�Y���:zJ^@������0Z_�;��ns��u
rf�X��$��s:c�r��qq<2�Z ��BFB4cxPb:�X���Mc�Q�����m3��Չ��QqF��4p���mr�s�xg��|���v��(�4^��.�p�!���