BZh91AY&SY䲘( <_�Px���g������`�{���� 7(�b5��	")�#h)����z��zM422Q�4�H���    h�101��&$�E4T� 3S ��F���4d���`F�b0L�`�!4�SL�Q���RzhO�=C  �i�I"��x A4$RIYP ��"��$U!'a2�����9��X� �$��e=n��}.��!�_�ǹ��Y����wwf�332�k�P�b͋�����<�g�*��OL�,�,����4�LP�B�=ffb�g�yd�z�=^���H�������)��,,�P� ��!1�8j[gi�s�����}-��q��(HȹU�yD�]:�J���+;L^Z=ښC��+uJ��'x�"P�ܪ͋�Bi���|�Or������E�~ݻ&��ZM�X�L{�\JR�)�4��0ޭ��.f��0L�����6����/߬@�E�g�38�m�;C����K�,0b1�	�'�������,���A��p��'�6�mǢ��Q�F��7�c$=H�I(����a�Ak�x
.��0'k#)pSV���^�-w���&[��"x�R���IY0oN\����ׄyL[׌��D#�K�ui��R0kH%�nq�Jӫ'iV�`��O)8���ۉ���2��`�P����8�D���TM(�nS*�]�/CC���ޝhiw��:���{�.�N��8ծ�AK�U��r,�� Ed���
��"�u����$1\�6Y�8W3�����Ȑ#6�|8&����鳿u�*�-�M�6U-��l��m��s�8�gz���w�"�V<GyY���i"�RSҷV�㽫\˻����������H �I�IUA��D��{����.��͆������O
�ρ�Q^9&g;
ss�!s{�y�2QTYJU�(�R���eE�Y����PX��(+�Z�)��7��9!��͵��E-Y����i���h�Ty�sKi<��e�z�J{���]�3�MkGru�(ַ�>�xSJ�����~����Vʌ:�q�\\�b��!��믫��c�i|~T�x$"�шG� 7�����Ue�D6��a���~�b~�c7�汭�=����;V��?�a�u؝G"�d u��Qa�ٗ^��X���k$B��[�##չks�r�	I�����L&�94Ni�J(,�b,V*"�v�Cn�z�7��5��o��p�w;<��Ai���Ҫ��ؚ��+s/ܨH7�=�gL;
�^��E���H���ҙ]zQ<h�~$Ã$"�l"�nTrb�R�R����fM��"*�3�f���H̴ψ�Q!̅w%oR���iP�F@��a�27�`oNB�mk���Ө;$�ni �8�G��z@h�S�!�IVGp]��yʻ�R6��CHF3#h�#԰�22bB���	�5�HE�94��E�?3��2q54�'��Aw���M;��]JC&Վ���F��9�V=i$A����u�j�3��\h9]�ʆͷH��v��D��:��&)N��x�3|��>H�!�B3��)ׅ��׆+������mb��<^"�f4u�x<xg$:������ ���37�]Ъ�IC���B.-�AKx�1p`T$�^Zy��,�"
K����\(��������R��g �J����!m✟:�Q�!b��"�C���3#��b���1��8��^SB�|��?���)�%��@