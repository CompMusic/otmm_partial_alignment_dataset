BZh91AY&SYBW4� ?_�Py���g������`^�_j�� �l��M�ʶHM�i�)�S�1�j=@茁��IM j     9�#� �&���0F&j""� h  �   ����4d��OQ�    �H�����4�3&���2�4Ѡ'e�٦��
�RV>� ���p�A@?D�I�>���I�B�P	����S�𧋮�|C�~��332�3���n�1�����3+/R�L��Ϟ�qVef�6%�58�V^�3���C�p]�(�u�y��a!17[��Т��uuw�{C�	Pp�=�l�y���b�t�L��Y�����WV�ц*��IX��JZݩZ�^dXe� EҾ��3��]�6�
K��Q��ݫ<	!8=�92�t�D`��9�ZV�!JҴ�Y�Yw��Bi�oW냣b��>f�f�g�s*au�T��r�oy5-��4H$R<�lݾ4��a��SF+hi��,P�E�����FQ�Zh�J&�e�жP�#���c�)�{�w+{����An`p3���ٴJ � �@$iJ#��{�![*M�@�]�-MX��L4#2�iai�$.�R�Ճ�D��"_���k��CK��/4�FE��Cn$��Գ}A���6�?�2���X�d�3o�ވ�>�n!�\���ad�kk�%PS*|Jx����j?;p��XueGw`��L�m�n���.t:�(�u��&V��B8jz��v�F�K_b�UV�Gm��m!^��!]���j��ŉ<���/*��!(��ː4ӛ���J�Vܙج��e2��IZ*����U�g��2Dۘⶴ62Çz��]�	W3+� Z�M�!�+�yW��Cjx�z.ӥ#�69�m��ؼd���04�"ʩ�P����e!�T����!l�H����T��{vt@��1�bzt���!�CD���ܥ嚐���8�:h�9y2���Έ��5��$�G��X��6X,��8�L���T�Rsks7��ę�1��IDQ_���	�����׀���$%R���m���*#X��,��5V��*"�Ab���5��PU�ᣆa)U ���Y63\`�hd��YtL�1j�],�Ʃ��.��mz�W��6	���t�:����[f�͇);�S��gϲ�����a��O�U(�k�� p�:u�2��>���-5T|���������	�>*��¨֗X���pXsF��9�tM��G^A!b�p�K7b�$.{R曎V�U;>�q{%Ɓ��༫�yH�̆{�F�����녝����ZJ���A!`s�4ٮ%F�L:�nL[%�d �E#֪b�Ŋi��R{P8P�,��]8�HE�--ċd$,D��A���be�5OAM�ӔL6�i���$����!wZB1�YQ�#�d��4	>����KlF��*�EJ߄5��"ֆD��X���H�6l�f.ʱ��td�P��!0֪��&ٔ�����`��e��$��`$/f+�M�!�V�`\$.�Z��0�R�4��� �mE���	I�����	���,�����5L�����6ɨ�a�PS����)oD�)�E"_��L�Fˤ�a`�{�N��W���+N$�Ff�����7�2���Č�]�$�w�KXƍZ5	XHHS=�k������ɈƊ6�sI��p�p�|�Xa��S-E�rK_Ή��+���U��(v�Q!T�7��3q�K}@h����H6樔-5ȓ		�T���~ ����4��1i9��%��(��Y"W��Q�AQ�����a�4Ҭ���vGͱ�$��#R-��]��BA	\�