BZh91AY&SY��S] c_�Px��g������`��q�{wb�  c�f�Km#�	"L� �54ɧ�e=5=O'�yF4��P���A�A2$R��h     �&MLL`��I���� 4��   hh"�ʞL��C�h h@@� JdF�&�CS4�  dODIE�FdD��(�h@=�=�$��i�Y���{X�.�'p����m��:F=:t����s��.�����ee����^fd��S� �R�[�o{��uN�Ig�s��w�+I��ݴ�!pܻR�f
�S�)�@�Ӌ�-�.���?�����w�g�n�hh�Dw��";*���(D�E�xw1*�4š.P���r�d�]�17^G9�Q�#\�I��ɫ�S�M��Ӕ�s�BDX�#%��4<v.�E[,�� Pfue�!2d�3�W����<*$���p�I�w@�]n�5���0�䙔�7-(�����7�vf�4�e�<���n��ǹ(T�c#��l2v���0�t'n��}("�h:!R%���RN$@�Q�7@���3"��t�Q�HiU���)8A.ڋ����[S���Jppu��#B$�4��U� ŴM<S�4��"x�D��(\8�w����m�>�΢�2�鮷�[�A�2�n
Ӈ��Vxe���JEC�5!�=Z9��,�聧SZ�8�1�on�[�����h�Q�SSAm��P�73TEl�2w���q����'cB@v�������۝n���"v,z~��X����D�h,WB*d�n:�<d�	��Z�9$5�+|�˹蚔�X�����k�R��i��Cs�Lnb����R꨸�ގ�)�V�f�>6����@�H���\.$Jۙi΃����X��rf�!;���i�N���DsI8F�!G����	湻�*@볍v�AUE��g��`����� (9T�Q`�YƆ��N(Ze�ii��MD��ˢ�n]���(�+�UT!��gLa��J�<���HF�9�����R:R,�iTR�dؔ�`))�R�64�T٠��%2d��J1Yi"��cB([N��ix�����P�f4go8�]�����n�
�C1S)������/�]_f����(���I��8���8޿L�L���S`���A����c)��Ғ�܈�����!�]@ƍ�����z�� �Kڒ���DY{J(;�4����<���_��9Z$.m��c3���p�^B� ;5��L}����%��T��C�V�[�6
\�RT����!��Uu�B���vEJBB���b����p�_<[����A
AV�Y���*�2,�&e��1B�Z���^�ɀu����Β����hy�,�&\v*�Z� n{6��%��P�Q]���^Z�������p� ��R4���9f�7�iU�l��|���
�6m~9�$l\��e�8��ռ�q��$+C[$��`I��� oKH{2�����g:gq��E��(�4�`"xx�B���йƚ� ��jq�M�3]Ȩ�L�B�HTڱ�d(����.@"��GY@���a��� ,��d�74M�5L�3fua�`\(��������y7�>�ur``���}��v�>Y/6q�؃��ݭ/��p�B��������斊�>@l �խ8ap�c��]�&N7t26'*b�%�w�&gg~w���t)�m7O�w-@��t���1�
��b���1!D�k��<-V�j��	Kk%8�t�M���aK���ߺI}�݌(*?�8��r�k��;S��I�.*:M�F�|(m�"wۯ��^B=��C]:j��)B�N?���)��r��