BZh91AY&SY��5N �߀Px��g������`�����@ �jr0��P���b��� ѥ<SC�d��F�i�	�J�      SSM��i�F�C&&�h4d4�a)�MSj�d�z���h�@ �A�5=G�sLL�4a0LM0	�C`F"@��A4e'��  4=4���?J�dE
� ���z��@������oP� q{+@6 
�xhq}y�O�
wq/s2s+2ffffe݋�����g��N�m�R�S�e��G2�uW3
��VI0��҂��]�G�!D8��C�VVt+W/M��j2�j�u�F���<�翓k4T%��'�YR������zO7GJQ&�^8�,e��q-p��2�߇��U�{1� H���iԹ/C�F�d���y�p�Fzj�Hx�U��MI�P��	WU�5�E��i��?Wz�g��Z�ٯ=�:�m����62e�vE˸ܚ*�[͜6��Ɇcz�ӆ�m�(*���p��f�Pc�BJX^��<l��f��⅃��|��D�x�2�� -�C�uo *����ԣ��*�#X6i�rpU�T�v ���Tn��Ɗ��Z�=�UZ�ĻA�!��R�0�z^3�Ǉ0��ā*�[Uy�+*�ClU�X�V�Q@�PV*�b����׉��Bw[v�n	DdN��I���7��-����1c`[L�^�!����<Bؠ��F"�9լT��E�\�)�a��i_�%�1��9;��L� ͌΀%.Jiu����Ő?����K�~��~�&�GƓ@��6"3!e����Ġ���^�vV"F��J�$'(���Y+z<d�����U�bRп-JoL2
{�(�-+�疛�Q|# e{����Y,���B8���R /���r��GZ���4?[�!� <ML���G 񓩳��	� "EK�����i��v�m�pj<:X:o��̡[z�5���a'l�<4��B��,CM�p.�qx�̨��	!�n���(�����&�m��8�c='Ȣ(�uUPh*�'7/My��G��SQ�jTݺ�-��H�֢�L��J ��inC{F���Lw���jd��T#Q�&�k&
��� ��]+c�uq�*.�`܊�W&� �*�(���95j��I���`��lhB �vX��I ��C�z��4�̛J�N��U\��de4Z��>Y�UT䰅tFyݑ��-�U�n�:�WG/��f���cF��� �y����PE� �%�"��� 8�g��Z��@�NI�@�{,ub�2��A� ����<�FM�h�63��� ɠ��i|�_j�w&6���Ղ��M��ڵM�J�Z�b�P��ݹV89Q�����ۧ'B�t%�AJ�J�w�	H�i�,�Pl9Ŝ�fL��)"��џ��2�J�$����,��kMmV̊�\��|��p�H,��@�_���I��;��2�JW�Na̢��ѶCEY�3��1,�i�'Q!�U��Ty��(48H�H��͘6华%Zg�S�`g��9?��:�&�}u�烷XY�L઱5���^ A4l7�#�$�I�+{���NE3]��c �$^�ơ�2�`��o�WFw�(���,x�0�*W�*���*���f����yQEf���&CLwx�hM .턐�k������Hu���LA���1�1��/�a��,A�Lh ˘�lb��� ���ӻ�`�	�Y<I�WI�R�� �U�*�m�&p�@J�p?+��l�r�����.?�5�Z�	^���b��%�*�DD���d��d��X$wxg�z�q�vPRV�AD���Wm�4����4	����,�j�����y�.i��cM���?�z���F5������!-��-�?�w$S�	{cT�