BZh91AY&SY��� �߀Px���g������P�f�`%g[�]�n�.�H��F&�4FI�4�M�jP��@�b@��@m   �  H��4h�'�G�����4h  �2b`b0#L1&L0D�Ц�)�S5S���  ���U	�(�� ^�Ef�ϼ����2H�QcH}�ZP�T� �_@�dz��5Ů����|��-���LC�U�q|�db�K;;�iLN�n��	Մ3$���)=u0͟I�0y ��؛6IO\\�� �#s˲e	�u���M��U�	 ,�`F��
vLEv�v��eLv۞l׃FW��%����<˘I���V<����V֓���z]�(U5T���%dzL���#]t_[/��쑙�ѝ脧�x��`i3�� 2�͝�h,��˥@��,PB�G@�(����$��i/d(&B:�S� ��R�n���@�q4(K�"�@�^0Uf�!g8W{������b�Zl�	�qg�8�s��p�c��VsIw2�k�x�Y��&���*��$̖�m~yl��밭)&�Y��mc^�T�����&�m�IA�o^$B]��*頪�&rZ�!ℿs%�P6B�ÇDBD�J��ivDJ��"��\��M�84Xa��CC�I�e��ɟ�:o���/]�t��7d���G��֛�9=�B��YןTr�M<�w[@�4(7��d�L���	�(h�TKl�h�����^�oN~j	 oh#��6�v����:������ve�%�1���nU��k.ݠsi�R��S׭��g����1h6
0?�D$�*{�T�w�����@՛\̅�ta���+e���m��S,�Zo�FI���I�`��dv��#22֋n��̝���2-���(T�F��47����%�:.�d�؟c)�B^���ָ-�4y�KL�i)�8�䆸�Tn��j���ޒ�!�?QV��H�K�a��DoUS�D�Q�8qP�M��iX	eW�I���S���P�e*1e�����Y}MQD���/���&�)M��#`cy�꿈��M%���M$aLRa�A�b	���6߉")\80�`��y��",LB�
�9$��Sd0��E�a���f�	�.�2�{��3R�5c�H>�WS8e�r �Z�5��-#nu�)bY���+�� ��\&��]�h�n��<x�F��C-@�����U��eQ�Pn��ύ�Z��j���}�p�Y�rz��9��%W,��9�a�#4��e/����%�S�u���PH�ɪ�a2K�7(�h>�C �/-���e��;J�a���\�&�Sm�ฃ_G�n���
�x�]��B@f�@