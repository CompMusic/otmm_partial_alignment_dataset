BZh91AY&SY@=� �߀Py��g������`_3�sp ���� �S	����FL��4���� =C#M4�4h�440j�� h sbh0�2d��`�i���!�JzHI2S�2mL����	������&L�20�&�db``$ L������S�O�T�hz�4S��=$��g�҄�@$%b<�	q����`%�!_(~a�4�E�rd��d UE����/g�k��0���Y��Y����wwv����Zkt���p�S���zP�t�Km@\�f;�\5u�4QB1W$-�2(���%��0g/A��s4q����Çձ�~E'!!.KBXr%��ژ���=�Ѩ!cz�%3��X e8U��G�u�\���Ӵ���%Ő���B$9V�*�)�3D!���_�LwH�")��9���X\.�/�hL���w�/5��QE��J�t�G1�s��Ûw&݇�4uXނ�6�e� >K����uOWK����/*E�B�Q.�"����*�n�E�c�C�jvnx���j!�`�C�e��#(sRThQn=b[�>�QE�B*�����0qL^�s��2���v`�SY�XA��B�R�6��C^��',�5/b�u�X oJ���Gڇ���N�Zs.zf/U�k�3�A%A���Q�f��R �lӍ1� �n\K��E�\f*�\R��u�z�I�"��E	��[�5\,V�n[d>�XGW�YP1V(K����fYp A��r�He<����*CX=td�Qb-���DH^����ꕷb��#`�i�}��=tp��Gh�Ւ`t�B����\t��Qb�<�m��v�:��Y�`��"�����su>��Sn����	E������SihPv4�m#����̫�(�!Z\E�!i���E��ֈ���e��kXm/2)!ɜCI�K�1t^s|���'�Յ@
q;��l=�kh�IG��a�}h�}{|*�t�f��/>���J��+?嶌R(�2�iɧ��z։]ںU/U�F���ڃ9w�G��kqHE��(�.%y���儃��1� ���!V>O���r�[�����^�kaaܿ�A����f���d���L��ٵ9�\�u���������޾:�09�[}�ˡ,ZR��ZEADk�!Vv��.�CI���w���Z��!�w�C���ޚΪ�"���b6a���VzD#�5���<�5�Z&yY�*&BC���H�m��Bw�1�9�F�]JV6��1�)����Wj��F�[�#R�!쐆ⶖ����;�]5-��fq�섑0�q� ѫ�\T�5Z�B<Mꗌ-K�4�[2���V��`9�r
��!M[�X���	#TQ핿%5[����a�3���Ί*Z�.(!��n�b2��	����!�����l��؏�m�_f������8�>���6�HE�����Q�B;B�3�ȧfm:��y�Y����ۚ�y��n;ͬ�F5��Z�faeD��QH���˫��ˤ�S,4��%���_�բ�5]71�u2Fk��u�����R�R�C�cF"�쬫�cqjB%$�A�Ls/l?�U+e�k�FuG �ϥ]���"�(H �g�