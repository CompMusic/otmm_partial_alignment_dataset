BZh91AY&SY^y4% �_�Px��g������`.�;缠 A�z�0��I�4LS�ɤ�m!�M hz �@	%5����  h �4���7�f�Ɂ �0��hh$�E<��� �A�  ��bdɣ	�bi�L#0		5<I�$�oMM�z�� �Dz� +)'�j P"���$c��%��b(o��NJw��jiA`�Qe<��?oS����dׯ�����wwwwy������uQ��`-���W)���<)��\�ڇB���i�����,'yW�*T;;�b��ʰ�H��8F�;14Q��D(
�H0��4(
JUز�J,����v\�U���T������
p�xI�fw�a��7^ȩ;��$����$!��^��g?�4��<G�Er��k���Mȝ�s��j�UV/Y�ōd�8/L�B���/��Ȏ�e�28�ބT����ճ@�9�$�����>���q�l�9�!��*0��6��廆F 
$B��@Bˉ�P�6�K�O�*+rwwT�<�PÖ���u�L�E[U��5B�y\��݂Ӱ]y�<XV�5b;%�E�|Ga.��~;��R3�6����HP�\]{u��
.p0�
 8V0��(Rl,�R2h�B	��j1�ЎN܊��|顯����RE�&I=t��ټ�0�(9�T읝�k���=#�k��3�*��Ԫ���44S�->)!��Q4��WWa�S�q^9���x��7���2�?�&�W������:�Tx.bE�q���v�'D����Ǟ��tي{QL�ẛ�\�Nm�'��/RChaM��=����ʺ�݋�y��_|��H �K�T����g�ޥ:��h��f�y�N4̺�T�Ql-�A(�١-�搜eJ����iZ
�T����ȪEE�SL��Z��M�<Y�2�fD���pH)��U�����"��=3ٙq��m5O�=��cdh�B���kθ�J˓�շl��e"�\Y�3;/�q����R�vo� m=�<�YٖS]f��`�B__<
&+]�"@�k{_R���;�%��e�t���m��+�|3���.1�_��o|�r�{����j� �R��oE��Մ��1��P�Q`����*�'M!g��X,�T�w(J���/jRސ���C����3V�θ�u�ѳ��gP����$�י�����.J�(�I����.*�L�4շi2ݪӴ�\���:s�*3�)6��ݻ%��=7/:TK�
A7x�#�|�~I�ۓ�JӒR�J����B7��]dR�&�w�v�0�K���Hŵ���	1`Y���

W-A#Ġ���	�T0��ovꂾK-J��d�(��U�λ�v��D�iJwo�n�T�ǫ�7�;�lڕ�x��i���Pm�I�q����`����Mj'0R�UQ��\�{����8R�C��d�̍��:����:z���'UT��$"���s̿=����9�qsH��erEbJ�3�\>1�2��LkL�p����qm���D�$Aќ+\[q�mL��5��[:㔢�4zQ��.�p� ��hJ