BZh91AY&SY��r �߀Px���g������`_{sw��w�} �7ϳn�D%C��(��O*~���f��C�=M4h4���!EC4hd`�h ��(��     j"�T�� �   ��dM2�?Q= ɠ=C@6�����"�55=O�5O��5���0M�'��$�A$���!{����I8$�e!����	!4 N�'��h� &����Wɋ�.Q�.Zg9�s���fff]����ffehk�P�ߩwu����[�fW�Yb������ZUfSL�A��m��$�{5r�ٕ��./0�2� ��m«í�x���e��`�N��WK�4��E���("��.L�,�p[`	1%8�\Z�c4�)�� �$� H�5i������^���ߡ�psË�fm(�&�&��C��Td
&���[RHi�7�O�r�mv�~b�]�g�<ً�L����,��6E�����JU��v�4�҉Ot�-*��,(��ix�<��9X1���ē��QM��7<�	WW [ҖF?��ʰ� #����E��T��AR�!!�HY IuE'����+��k!wU[)w/����"��¾�H1J����hjlf
3�&��v֫� U�a�����u)�EЧpFol��خ�5�R�ʔ;���̡�F���M��\���oZ"Z Ҹv���K�V��Qd���Q�Hp�0�ځ[�WW�-�!q��?moa���CZ�_Y �r��BI���_�U뗑�l'{�!G����cEE�r)-<ۜ�-�%
aoL]R�Z�����*7[�F�h68i�7,��]�h4"�����:�S�E\T��S�鎎BT,n��FDf<XN6M<���[�0U��� �MK�q�w��H�b�S���:���0��@���(�j\�V��-x��1����Cw-KX��wA�cy�m�8n�k�!��R?΀�Q������"�.� �,�k\5�Z�hM��4�U))Wz��q�-�U��S)���M�WMȱEb(6T�,�a��هi���P�$ڇ
�;��2�a�5V�k@�H&�1T�������'Eyw�̱{YlHf�kFh�%K��� ��E4��
�=V����/e���7I#)L�ya�������	_C�K�\2|�G� 8	[OF��-;h
q�6y�I$q��������`����ښI\�����54J�\t�A��SM��;Dz�(�`����'���ow�3���Gz�z��kTm�,��bB��J�"+`a��3���\�Y�e)�k��d���_i�iU$�CcB!��X�KlMS�O�əc�oN+FΨx��YP�]$�n"����[ғ���}점`
�
��}��_b��R>�JYZ:�QV�R�m��Ǭ��j�e��AQf�¸�l)яu*�*Xc�xh�-�'m4�ke�|�$�O��!H�֒G]��F�ͳDCF��TnlI#��_pђF�р,�F���A(�6!,����"1��H����?HSA�uEFb�z�^�"��Y�ܪI�X����#rI�(���B4)0��!ٙ{\X�A��!�X��|���y	un()P ���1�SڍI$y�RH��|�x������e�*�m�&s�@8Rp<�\���J�6I��+�q�ܶ(-Ԯ�T<s�I0�A�M���e�C˞4�t�Ť�g\$�Y,��R߃�V& �)��;w,Z��$y>k�֬��n�p Ru��MG�qU�0�ƿ��3��zi`��7! h�rE8P���r