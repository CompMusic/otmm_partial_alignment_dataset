BZh91AY&SYGz�u �߀Px��g������`�{q�F$ |��[I-4��H�hL�5��Lڦ�F�CF@Ѡ	&�4      i��&�&	��0`��$�A(ԏ�M��� �6HЍM&�4�  � h"���6���S�zO)�� ��
�n�D�"�AB� ���K�L$U��$#)5��y�I$�@^W'S�L@V�v�}�8��m��[m�Yd�������������˦�������9��WuOH0m�����'�+�C��[R"i�
���ۀjꦑ��� ��ⲑ%8�y��u=.Y�xz���Vh�_3�7c�* �>؄�%B�$2�;ej0�qr[wP�re���LNo��rB�vP���E�:b�T�>�ak06c�B�D�̢Xh��3����F�D�!8(�s��vI�"�>�d�;��ƧW.��_k���3YL-��WV�믌u��;���eaK�)7en�x���x��@h��l�KƹV
=�S5��T[t&C2���F�Ff.!�^Ln�t =����@�Cf��h@*%�tа�IL�w��y��i)�cVK)��(@���ax*���˕ntK����x���h6�\G�nS3��X/2�ʑl��C(m�<��*���
YB�����!eFD1�lW�@3�n�����;��$N�I�\���
�O9(��lJ:0P��LU���D�!T--c�N�����fp���ku!�Jज�p�s)�Ts:]���U�F�ȴay; ��H�� M��\ʾ&�%h9;����E0�bD��p�<���?�[ho-a]�/^4����_��P� ۉ7pY5i�7a����	��U���N VV%�W6�H�"N��{��ؒ�0�L`b_9�A7�WO� ��nLqj^aЬ���C���������a��2h��e
�
|=�7Y��N�=��U�[�]U��uXMъb���=q�j��;�Š�$-Ep�P��e��|�
��ˑA�HE�޳�|�DQ^j���	Տ~y
c�Vi��C�!�5�t|�
g4\j��RɄ-��Qi�*6�j�(�o�T�2�TE"�x��rL2�ɻ���e��)�m[h�m�kL�g�ɆF�ܯ�6$��ڲ.�������+��|���\��r���H�^B������q���.%0kQz��4Fa�`�d�N`fL L�q��ߺD�C
 �E�x �ɿD�D
�$<����t�<��M�VЗ��?��B��}�f}t 溤������������ �Ĕ���B�:���|��Ow���W��ѾD�%�\tM�HNG�f�Lsr�	I�۵|S\��aP�:4�LhX)FA`*������R����o��+Y��4L!�?<��-U�$(P��6�o�ֵ^�5����մlĨ��f��8��;J&k:�̲}�p�c� �:	e�&�����\gI�X7ԭ#o��Ȧ��p��x����s8��f���f��{&<���V}��/%��u�uk�kw9�FXE[j��c�N��$s�cjuʏ#k��BcS��� [�O<DIpR���!�i L�T	�Gl�
MR=D�EU! �?z�9 ɹsI�i�a���&f�&�(j���+�kGbHZo(A����P�����X���p5���e�0�È� ���C��Kf�ld�hM̐3չ5*�-�$)�������7y�WoAxy+Y"��Г4Ѐr�ny˔.jl33���"��R�Q�3�v��.�y��qw�H �$"���#�$�)�w�PX�B�r�	ҋp�JG>���0���P��+t!�Q׀�;���� ���@x�.m᚝L���5�q����Dr�e/[�rE8P�Gz�u