BZh91AY&SYZ�  �_�Px���g������`����|�  @�{j�!�U�$��l&�=OQ�ЏS@=@4�M� I(��h�@����2b`b0#L1&L0f�(P � �@   T�Q��L�M=�h�   i��H�B	�=��S�)�ڞ�������,�U�Gv �*�
��a����d�6�$�0����� �e�6Ds�r|u�'J�{{���1�c�fe��`�����˶ww��1�j�P���w#�K��j�&	i� �R���`��E
	Y,�mS��JZ����І*�D���חٿ����
k0d�U�xi�#Yr�6Ԇ���4�(hml1�ZR�<еAIQ�f*��i�e���f�A����V̚QM�P����@UL ��Y���	2d�g���bs��7TR��ɒ��h�I�2��s�\�d�0�%�*��*�TY�OK�q�H���1$�,!f,l�Ue	���4#���k��*N�:�j@�����r�x9[ܫԅ<P8��I.��L�� ��>��HʊHI$�-�H��Q@�(��ZL�:�1أ���S&b��R�FEƫ�)2�3&�V���Z]š�.�ZNR޿IM$IK�L!��3e�f�Qy�	�/X��H �3Ų���cR8�o�
��p7���#�^ۿ;� �3_��vt qT	(�����AN ��V6n��dT3<;.�F�u���$t7�F	E --� � p�N|�O\^sY�9��u�j��h�kw8�Q����ʘ�,i�Cs�݈�Gl�j�
f񜍕��Vۗ��i��6p(�K�(TK�l��/(�����xax��n��9.ʺ��-�u�H�d5+>ukqA�׾�����!����tqD�=���(�nvP�_q5�0�M�����,?m,�����ƕgE�6��+�!u�9��#j	J��ޖ�P����� ,�YHq7�Ja�t����
���kq�l��� @r@ Hm7\�^��j5�����K5M������� �0`��v���n�#t�#���v�jɲ�F�BD�7c���&� H<R�) �DI5��	 �A��(�  Y%���y�)��r���6��.֭kBM�&bvT:�����x���>{qoP+�{Z?_̏(JևZr{a49����
iR�j��w�u��VF�6wI�i�3�]�l�]ŷ ��UN��A軪-I\ Cb" p-�<:��z�<S��@��X��мF1� �`�b�!*.u� ��>�m��E.�3h./�tב-�)>ˮ�����ʮd'�t�=
1�F�K�.�ϙ��F��_�	lɥpcm m�La�����h*��D9���vL��|j�p�4k��I�Ҩ���B���pڙϩa���P6��6�Ġ_�eBB���!�ܓ?z麩�!*p)@�%pm��7r��(鼄�_��$��JE�]ӆ�&E�:I��X�:���	�гJ�{$$�cUx����n��:Yj�88G1k$ <�!.�+���K�!��
�C�[!	y+�3H�B[BY��c#1���u�&X�ζ@J���PFUV
����	�d,UY�f���#)ڌ�w*!&KVd/i%b.��:�̢b�0�v��Wg<eb؃���k9���8�Ak�of[�D�BBX� 4Lb��G	h��_��f8b���=VZ�V�ܤ���£��ٞ��C֥&�4����,�d�Wa�84�S��sS�q	TǌDMD�@g��Qp�i��``�%���N��~��1��L���m�΀}�vC��c�D�6��[����S�3��ʦ��a�'g���%p)C�TM�rE8P�Z� 