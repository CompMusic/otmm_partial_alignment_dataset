BZh91AY&SYK\^� !߀Px��g������`	-׺�� �+6�b���a$)�MFS2�����OSz�G��46�#mQ�4�)R1�  A�L ���Q4P i�@ � $҂JyPz�C@dр&L� E$H�6�OQ�i���h  �M	=���4�1=L@@�6��t�J�x�b"@�}G���$"(T� }�;�܂#$/Sk��H	��F\�\[m񻻔�)p���Y������������Y�����Y���:�H'XP�����"��<����06�d(�0n 2��-C����OI��*��u�*�
c���]g�Lፀ[K�ݖ2�od�o=su"a1f��S��a�E��1���u����7&:���XQ��ai$	3��5����;f{YS
�u����V���j�iL|��%��r1�v�
�X��\W�����k=on��c��]�7L��z�c����`�/&Q��Z݈rۜe��eC@`Ӽ�ve6!��6W�LB��0��>I�������86��e{
�#�����+T�U6�U�uq�j�D'�ns6P�A!dt6$���Қ�a�a�a�P�(�z\��TGc���tz;�nˉ��5�8�7�r<T釕9O�d��V^{���z��x��P���.Z�Z�KӔ@J��aH 3��0CPe(cer]�a@nC,��I�TkT��f�-D�X��Yg��̬ԕ_MtW.�91k��A�� c¿,�.���P��	 �@�K���ʐ4���|����1�5ý`*��"8$N1r��d��:��]��4�pDT�a� ɉq��q�n �ӫ9=+�В�/��m��A���:8:�*V ���6-`l[8�Z�TTO�=h���JZ*�s 2�8�_JrB�Rya�20�R���n��yC,�l��&j,8�g���>�L#�*�NYV���'5���QU9�"��ض7@LS����aֈZPO+Q�)��4V>']�^(�����[����_	~�Tv:�Ljo�^�����ZeU���5`v�G
ؖ���R�rx�;+<��>7	�m2h�^R4�� б��e�+���∼�ǨH �^�TPa$h����x��6��]���M�В7c��b�B�AA�(<�qyVE
����U�wU��b�D<hi&y]+$7��e���7jwN���%D�hadm�vZ��%�G�ѭ�0$�Q��}2{���i�����k��/|?�->����a�P1���̻����T�h�-y�zy�7�����s7i�YC��^��a-��|^���O�m�ܼ��	��! [D%'p�٬��A�
=��Q��%�z��v�f��ݡt���d�O�V/�A��̘��D��Pk�w�Ⱦk�|����	
��!��n��J���&���K��	-�fC4ߓD�"�p�M�a�	6,
��*�R �2�O�����7hp��.�^2N�Sslȋ`W�F(�%}���2�R��}H5gg�1���P�Q5�YNH+�I$�G��/X�2Yi�A��_����G9l
O-�Cw��N�I�3�LXXr�g��[;�J[��u�2��&5��=븻��mr�
�1��3�o��N�x7��7�<:u$�P���� �G��
�u�T"j�^`4����@�Y�߸D�ҋ�]��n�T�fPW�����v����bBD�����ڨI=6fC�' ��s��+-�zb����CT�E�)#��Ê3�}4�����f�� ��/%���`.56ʥ(�i`�FP��H�&,!�h�ad�Ӱ��!Fn*r&�W�/p���/��1�ϐe' �B_#$.���U����;��uN*�6����F�*⭧J�5'jWe%5t;�<]U��B"��ih@�Õ�Z'��A��-W
L��? ����L����T����\&qkM�g��fJ�Y�J���̎�jV�I��|Y�s~�%�
Q
����)�Z��p