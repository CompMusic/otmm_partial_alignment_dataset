BZh91AY&SY�Y� �_�Py���g������`	�������Z )���Ӷ��κ�I !�4��Si䚇�M�4z���=M����a6��� �     i�BR�� 0�4� &�$Hڦ�M�h�     ED)�z�&���� � "Dș&����M4�� �2��F��RTU'U
̀� 2���i"�B2��c���@cx\�X6
D�r�8><�#n��%oo�%m4BdITD$�I&�̒I$�I$�P��Ç����As49
Q�&�!L�/n���~�b��̣py�6�M����������a:vL��E ��煾[h��a��o$Lik�M�����|Ș^`�iw�B���lui[S.��M.��-�Q�%p�V��l��$T�� H�D�oX��#�{�^kY疰�Fi�G�Vq�'�Eo��)1��jP(�%m�*�݅�BM4��u���Nckjce�j�WߖR	�_|��5m[�F�a��l����f�5[�c���	5M�q�"6�`/�n�A���DP�s���(	k�J�q&
�#
HDXE�zV%��R� �u$`�"�p}�+"��X)�%�
LC-���t�<
�tC����i�Y�\�I$!�I��)�	��;xEjQ.��)a{����	����@�8�v��Y���Y2�Y�D�Aze��f=��	N�Ӹ��h����Ա���H��3�����VI���y�*{x�8GZD�`7Z���@4A`h}��\�F�;���Ӹ��J�M�B��l����)h�ˀ�1�����I�qb����/����A�����������:<�rF�T����L:!C�C;�A+4IN�\E�#�p�M����k���[{��-��	^QᎶ91ǰ�UC�H-ZJ���8{�W8A��������9DY�g`bb$�$�
ֶ�Im;9P�uqV"�fr��b���J�a�}[�� �M����(軾�m��mӣav���7]��2]8�O;�&�t�^K�h���b�xj
{��q��^�Ns/Sx ���4��>����S�gĿB���^�l �f`V{���T��zt��H>Ƣ(����24O��=�Xr�%�{sa�������=䠬ࢵ+Z�ckDie�o�8�W*(��y8�d�7��L�Qb�L����ɼ,� �x��%M"�k6Ӌ1�#�*�䇕8g�z����w�蝌�PNl귮.�{�4���K8aN*�0w{K������hrNOmq���YᏥ�)�D�ߋ��r�U���7�^��HK�[���������0t��:^��e"88*�w�ZeH�4�0]d�C�˝}F4[ <��!,��ݜ�sc�rƾ��Z��t29|����L��嶥��l^���	6Q9UZ��%���M�ϋގ+�ۢ{� �s%9DA`��B�
E�PY6�L� �i��eY9��zd�����2��%������������W�U���7423C��W��t-������H\�ⴥ3ʮ9E0�d��l���F�u���Ҡ7-�&����
�3�w�����Z�|K,�&<�[�t��WQ^��V����$$�^i������f6YW&�h���hi 8�%�ڼ@4j�_TDA/�LИ�:����g��YS@��)��j��,0�,�H	�Y5������0p������~ukd,������������I3K�`��6�5�'�d]j�J�u\#qU����J��l"A�Y{��Pm]ٍ�1��y��r��&X���� mɆ�܍��@BQ><	g����;tQf@��<�mb��<^"�f4z��hs�0�}��XB�L����pOj��!)Tז��E/'U�"� ��it�n.b�/��y �Z�)m���0�!/T����~
�A�����r|��zT�E�ժ!�)rO35�T�y3��f��0B��h�_�.�p�!D�( 