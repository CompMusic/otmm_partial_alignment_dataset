BZh91AY&SY��o= �߀Px���g������`	_0�x�J  @{�U�P�$�4�i�����4�6�@�x��� I%�� � @ )O@�6�#!����b#)�L�@h��F� � �9�&& &#4���d�#JM�=M5Oi���2�z�?T��-����` �P])�Q��S������?�'�=�UCA<�h@��)����]���x�5S�GǙ���wkw�wWp�/333/ffe�ت����7o���A�N��9���Ұ�*L���`2��=ئ�c$�b������GL�XB�y���� Q=DX�5UWB�2!�=j�*i��'��m$�
2}pI,۷����r�ښ�íP�i]�#>���	楩�	�K�&b��q��խYBe�2P��O'��L�^��j��x����+f�vu��\��},��3B�[.^S�%�rNu��7��$zIn��/.���&��w�A���a�e7�I���r�˧�ޗQу&Y�h��(	�+[L�f�X�uó�UD���[\��)��hh|�Y��WK�Rd]�qy,u`)z���h�x��Z�/ 1��d�nt8e��
��bf�yV����K	�`p�5s��4vw�1�fX�3N��=7������t��9Lύ(���$�󑣺��L�v���i�*�p�K¯O~�VMnar�1�O0�.R�[Q���m�0������I���5h53+�pD�*s�;�u���pOR#k,�2��RX�v,K���vZ���#W�e�7;�Z�J�T�fY�t�X{|뎶�TZ��mAsJCZ�)x5�5i�
4ݭ�dIQȘ�%�r�`�]�ٗ:���:��6Rސ�ȖلG����_��
��1<	3�|��-�)ԣ�0`��.��l��6Ր��3�Ԫ�n"
C��C�T˙���x8���̼����\���V���J�՜���ጵ��dA�q ]��8b�n6pf��qẖ��]��Cw'�6�;v�VUn�����]�w��R�h�=���A�;B�3��P�,��v���fn�V\�`@�h�$�[ܜz�e^·h�l��Om۠ѯ��S�!�%��"ªv��2b�½�#N��͈�Q�rw����hy�ҡ�	�-$��๽��hPy��*�^6�TB�*����n�_��;�"��*�TPB��xew�U��ɢ��}��T�ڃJ�B���B�Ҋ��Јܪ��1�
�(�KQ �-M�=�Q�*D�8�(g!�Q� �Eޱ3�7�wU�$i�]���k*��kBu{��u�J���HD.#7�q0���Qc2��_�pA0�2^�8&��42�dGJx�c��7n�7rz��xJ�9�Nf��������z�B��z�PD {�S���M�3<-��3��:YD ��Zn�Rn�<zG՟Cw���v���Ӽ���K~��TO (����V���G������,����}1�O0��4���K��u��s)#�"F	�4�I��
���H)�:��"�m:��4��z���PYEk�N�[����n�̐�@��C�D7�r/Ό�S���>�L���Z�^�r#���b7��Q��C�P�I`ݗ�&/*��QYe�fXƙ�)^�,W2B¶�F��?^�vR��=�)�v��:�*8�{_���ȳJF�]׈�{���e�u�L"�i�D��B�I��6�r�	y��S��ˆ�Beq(R�� �΍F����1��_E횲��h*"����bt��S���)�<���%�o��\h��-Cz�`K��zG�Dk��N֊!�9B_����"ဈKX���w���c��<5jL$eS���.�'���:p��^|�� h�\e���&9`"&D��<�� �;�dc[�!ĭ.��&	"�i�-�l�zB4؃YC#8�LMe֕� u�_c�![0~˦���0���#�����h�jFL��H�
;��