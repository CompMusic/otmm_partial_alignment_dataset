BZh91AY&SYX�� �߀Px���������`_}�����t ⬆T��S�$�F��CЦ��jb6�Md#i� �� #@2 ��2��2b`b0#L1&L0f�&����2��   ңj�M2 	���h"Bi6��ѡ'�=4�i�FCL�	��`��� �IQ	@�}}ė٨hm�@	�4�N��EI��&�PIU�w�����?u{]��vg��e���ݜ���̻�����̭������"1Gh�w�c��;!�=��UEE8jQ�X�A{כwmZ�Z�Q��`�V��w��L�^��A�D�H�>��!]T�$�b�H�$��2�p�q$d�rp7HD�&�'�(U��5_󈄄	Qbz�VM������>���>z���dB��qq���\E�I"xQ)�<�V�i$2d�5��ִ�&0g�ISm�`�^��KvncK��D-�Ɩ��^B�I*E�%ܔ�F��26�����؎A�^���B�2R�2�1Fc�rY��h���,���P�>v<"�/1�P`ch'>i4�p∖�f��Ű������Gb(Ƀ�*!w(�YʦV1�	B�i���jbݲc�V)OF�(pm�fJ��ɡ8F�� +4�P[nh����1:{7N�6\�*�lUEC0um8p�(4HGwl�BQ�b4B*�p&��6Qi�3��5-�/���8��xJ���EP(��]5�]'%��������up��Ln�e���P�N�P�/Aj�+q��-/Xsozu�����3�Q�)����B�X�w�`ƹ*V�1v��q@��n��H��`����9m+Tn��Z�;�*V�Am��u\t��m`�s�s��]:Ѝ(��"NuDq�'��P�WF��v��B�N�	�W)7 6�&<kr6)"C�qm=�Y�8Y�O��&�˘�]L�6�^�H�4�v�h 		$ȅ���}�5��s�V�F�U$�����T�]%dR�`���R ��f�,�MtD����Hƒ������"�`�Q%B�T�ؕ�Ye�g`N!4ҫ�_{\�4Q٢����؄3���>-_S�Z]򮝙kڠ���5w��=#t�Z>i��|�_�ۿ�P��52t`x�;,�	zS=z߻b��Ƨ��n���j�Xr�����I٠im X��_I	$}5��>Iό�Ы��=/"��T�E�W��� �`�Z�K�kL�E[��o�F��c*��S�$x=RS]�T��'RW��}W�;e��3��F�\͋�n�f)b]jk������N���HHHm�c���I:P\9�8�*�Ͽ*q�T%dv���iQ$�"!���Q/Q�WŻ$��~diX��=��6dT���H*�GuHE8�?�lK��5֊	 S�8"<36�qǡ]u�8|B0�$*�N�u�۟A"W/TN%%Gp�ծ���B�$��3 &=Eο|��lK^��h�k��z�%Ñ��!<ՂI��(���I��gqJ4�)$��H�BZX�dkm�p`a�A#��KQ��H(�<4̘�+�mc���b�)'(j��Z�
�C���u(C&��E���h�$��rh=�u�
o���:�_&p�խ!��5E�s����8(���<g}@�� �ŏH�I#�Q$��>bZ2Pmې2hAPl�Z�3A&1�p3ޙ�6~��_�֕;�v��w
z�c,S(A9�m�H��Q++&��P$�]}18���Hq����e�I!���fa0�M���1�K�ZI.)�l�P�H�Hݮ���G�ܩVV��k���xPK0W҂ߠ��)����