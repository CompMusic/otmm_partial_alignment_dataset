BZh91AY&SYa&f� �߀Px���g������`1����  `�rb�BIh&��LКe� dz��ښ45% 4��  �  sFLL LFi�#ɀF	4�"SF�=LF@�i�h�&�)�)�&CC#M   2�D�	�4�4�M��h h4�ot�$ �$�� !	�:�����B�$���ID�I \1;,��*��z����/wx��}l�e��UV]�fffffd�*Ъ�����������*�~��g[�.�,�a�̘u*U�AuR�+U����邏I�� H ���{,���=N&P���,�0�ec)d��fU��C��x͑)�m�&�-xX��٧(�Ee�g�Լ�KZ��t�R���؎끅�BIĒh2�	Mۣ�I&L�^����:�R�Sly�{Gc���}�r�G���ZӪ\�i���n�˚sX�T�"Y�h��6��GT����M����W.mq�{�$�5�8�|1����$Le��)�׈lxD�"5����Ɛ��(U7b��%�
zfq�,b�+���0� 
!�y�C�j�M�7�ãuT���,�XL:ŇBp�]�d0Q��]Z���w��S+skQ���T�؆H��$,�v3�
3��pY:��D5��-����85�%ЊUշ���qS9U��vs�@T���*��m�p.�I���	ڇG����Yr/h2���:��1�i���2̲���т�/¤R�,0�XY~\[���8es��Њ.��Ɯ�m��q8W��ru��%P/;#^O+\�,T�X�)�$;҅eĹ`5�����H�#�d- U�Eg�YP�YTӰB��Y�E��-���-��h�R�h�h[���,@��OP�J/L�Pt@b�Ȑ^�;��۵s��]��G^�V�$��j�`M�X\��ý
kmja�ŀ
x�7[�DGZT�:7�c�BCI����w�����1&�jz<�[PY����єAa��o�é:��>L�V���(r%������pn ���28m�+�
�c~F�4�PA�|��<K���l�I#U�v\���iQ�[Mf"�*�����"#l��@�n�z��R,X��.�<*���4�l�&�E �J�"I��l�DkD�'��zw���f��z���L� �A�uo-�;�&�B{)ے��{�����HI�9Ke����'SI�Ĕ���]њ�F�p�=������1Ϲ�[�D� �X� 2Y�ȩZl���ׇ����w���$�x��Y�Yw�pK7��y���)����(RR8�#�.+��)q�n;x�_��L���J	%��F��D��R�i��Vh�a�e@�PEV,�b��H,��
 ���E�X*�'a@��k,Ԅ��$�:L�_T���2���y�l�aOC�^��py;��!�)�I{&@�����Q�˓�h�$��U%�M��%��)��	L
��j+�h�c;�Z!��jq$���I&*z��7Mc���}+5:G8�1���$r�%�o�\e
�����XI.ü�+�a�Y�� ��`�Z�͂1�S6]����\I�������2�]5'�,��QYM:-n�bI2���xs� �X�H��l,�?۱��n��u#h���?�C>��H�5=��b��W� ����`�[BbIR���Wm�����͎(�i�6p�p۪3�8�3\'٫/��Ȧ��v�S��cQ$�XxW��!�#�Y`�nː�v,��]���Z*m׀W��b� h�ذ� ,P��� � 9j���3%�]�,��c]oT�6�D������|���H�
$�ڀ