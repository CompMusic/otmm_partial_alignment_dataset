BZh91AY&SY l�4 �_�Px��g������`�{w�;�ަ�T`<�12f���Bi=��F���h��di��4� H�=@      5=4JCM4 24  �@��A&��A�<MMh��&��mM�12dф�14�&�Q�jm	�d�4�hЁ��4�f����OwD�"�D@#��K�K�U��$#)��x˒I5C��̀����376�p׳n���JR|�32s3332�s33"��UVE�h.A��.�ݠ���_d5���hr��.�U2�Hu3.���]T�2Q#�*X+���hK��w��َkj�{����c��{w͌s��m�8�I�J��<�^Y<(b�.8�j.�/i,�"������8�HC<($"�ή�uʂ���MHt�)������/*a0�7����#EGJ|2z1���δ�4�W1��~\�=Z:z*i��XQ	��tRs4-6�t��v�z(�+�cE���M[\WTD	���!�f�9110�0񇚸���a����߶�O�|�þ���3�����\�/9�iNY­��tF*3�2�a��d֞�UT!^;K��Cdƕ
@�k���.�IY+M�T����f[�Ja���Z����W�;��qN�<��p��F�4!Զ`hQ�0�	l]���b���
������DE��K"�C��n�	�uc�|�f�$�V]���ɾ��b"A!T,�J���q=��=�_͛�n4Jऌ�qk�L�c�nH�á]ti�F��N�Ь$���+�̫��:AZV�^���E����}xUȚ�s�Kf�n�a]���S��+\�΅2�R�^��v�a���(�e4.*�I	�2D�k�U"ߴ�bw3��&x�]���i�M~���E/�	�#�Y³X��)���0E�h�l���Z��KiP���+�X��,�c��UQ9#����nV���R&��Q4.��K4���-	"��$���W|����+,@�[8%�&��')�j"��UT$hN{���)�;,�S�c|T����6��Х�2͘")ޗIeJ�DP��PղAVD�����)Qb�E��`lZIvB�3i.���,J�h�Y�t��T,4C��᝘�0�a���8��jͫ��x������^l��P>���go}'��r�'➠����y���RT�5Qu?=�ϐr�O~�([Ҟ���U�Եi�g����{W�ԙ��C��"C��?&Ԧi�:ԙ�j��wA$+����[�9��G���0<�v�� ��:O!������5�AR�L�p{?H����-�X�yK[[^��:�;y�@R������'��D)�F ��,Pb�)'r���k)�^��hh!��8�Z�?FY�{����a���&�(�k��2��@��M�P�`��t�Q3��\�O�f�0�`ym��Y����v�s`�7��"�Q� )�"F����b���Y��zC]Κ�KE�ZRB�-`a��Z�x�vZ?�z�K>>`��@�|"�ǉQ����!8p4�I�\�A�Q�:[�!4��J�EI�D������d(�� �Z,���,B�l��r�EU2XOUM�A�Yi��%�����s7�h�K�&�GV ���j����Ǔ# V`>����`{bHu�(~�sV[���..�<�r��blN*��[�8aK�$.\RB��y��Y[�?M��P�ͬ�V+y����6�C����0�Q�W��� n��l������)]omE�0�gBY���>�q��k�mEq����I	����t�\,���t �~%��stBU%�ۜ� ��*���C�������փ�!�D�o��#���i��.�p�  �lh