BZh91AY&SY��� �_�Px��g������`	�z���  @{�I�H��I	@#FM4hFS�zMOQ�M42� I�  �   S�E4�z��A�  1�&��!I��6��  �C@sLL�4a0LM0	�C`F"�$���И��G��P����L�@ �$�\HFI$�~����M2(�0��y1���m @�4���NX6���-o�v>ޭ~���ka�m���̉f�ɜ9��wWv��w�����wwwwy���˨P����<=v�t�In��M2���R^bL9%H�w���4�X���`��e\�16���e��	8vH>eQ�ŤiZ>Mɡ9�Z�Yfu�ϼ3\I�͘a�k�a�+��SD��D2h!�52=NK׸9_��
��:@�@���C�Z�]�Λ˖�<,�孭Q���&(k'��Նcr�X@X�8!;�u�g�@A���3�������}�K~����j�{9q���,�1ww.
����	��l�`ݞV���il�����Gb@Sx�j�EE�A!|�\�7E_8n���R��f�4z��M�[Wb�sR�F�к�Y9^y�yo;ϡ�lɊ撐�q%Iч)3�1QwID'm���w�oZd6�y u3K�^�8Ղ�ҒU��o�:������e+�p�Y�w`ݝ��$�+Šቾ�Ǆ-,��@B�P!�fib/s1�D>�2�&��壉��u/&Ж~_*2��1����w��$�	�@W��O������#%C��X�dX+��+�3�oyӲ��� �dqj�Џ��8˧7&�0����^����YJ������d������A`8M��ܪ���L�����7Z\��-1��,�fn�2*9���6��;G�CN�G���n��ݓ�Wl��NC0*�á|�2����3YK�\��V��8a'�ƈ}QOAuh0Ze�:�p��^@�٘�|ZV:�6�K�y��(�|=�L�E�^7�8#�|K�)���	!�NRi��2Z=\�ͨw�*XF� 
K4���'P<K�|��<n/���j{�"
��w�Q��]�q�0�
;d��˜��)-�{��<,�n�͞wo�r���d3U5l^M�H��Pj1�G#�F]��Xz�L�E�# D�����+{�4����4��^ܧț��noq7jj՗�s-�V#Xڂ�ʫm����yZ(��J��g��h�bd.QU��g,15��֍��q*Ky+�1�w�n�bѨ�Ԭ����vwkhi�a��&>[�HM�l��0�9a_u9�
&����.���}�?����_/(:��t7�T�J���)���+R@�?�$7a�uSd�eR@P�ݪ�Pb)���O�ؗ� �|I�=$�8�g>��Ve��C�)�Sh�$;�G"�w�<�-��1 Oh��G%�j������(��'�Kʗ૛2��R�91�����_u!<�rq�++iq t��n�;��,&W���m�;�)xYܕF"�b�F*�TUb1!�`i�S�q��8�.ʨ�������h4` 4���Ǭ̧�bk]J��ڸ%h��[�� ��:	��?�IE�<��W�(^�v���>)�4�'���Ġ������Ҩ~RU����.��PI�D�!��Ӂ9>�^Bc�4G�#v��C"�S�^����� �j��8�q��u4���&���vI	M� ��])4^k!A�`�Gq��=
�(ѨŤs�ƐQ�8͵&~X��ĐB�x��vW����H�(pDCl@�*AY��;�S�N]ڇ�Ի��y�f� S�^���=#8�6݁*Gn�K@A��?�e����X$o,�"��c�]�b&q�7��}K:H�	p4����� {C Q�q0������Zuµ�ͦ�}{H%���n�a٪+b���6wF�F�`�l�Z��L
R�3�� LD7��E;/H�V�c���ۯ3U�z1 A��	MQ�����yK�4�?���d�M"� b�w�O}le) f�� ��i�#h�4���&לm�3�@m`�/:�ן�.�p�!���>