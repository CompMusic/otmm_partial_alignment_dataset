BZh91AY&SY�! g_�Px��g������`��]�� t�H֎�$��H�i�I�=fP�щ�h"*=&�&� z�`� ��&MLL`��f�j$H4ѣL�  �&MLL`��H��O�F�Sڙ4i�   �T@/�8� A@ HHN ��^L�m�%�!C��>�p�]�!C�2�w
Yk�jl����ǩ��MuU"R������������Ǻ���.�B����0jݥ�����V%CL�g�Z��u��ҹM(]��CvL�+�`bxX�������),	``�羴��f���ђċ��c9�*(,$KX�g8���tv�I�����V�+��R�nuީ;��>E�Yp�9)�ɤl�hv�]8��i�7�}]+�I6+z�um�Vn�Um3�UQF�
�`�Zv�*���*�T��
��5=�bGdm5۸��U�*[|(l�0b6X-���t�S�� wH���z�3���WE��HKc(�L�J�!<Ġ��H��>��bʁ�jT;:*$���>�H�R}(�3V�|�v����Aa�CK+��U�.�6a#�i `L;P7��KR:2$],�5���g����N�Uq
�fX0R�29�.ǃ�>6`q:�a-@ʱW;SN�K�`��A
��S2�%v,*To����A����7�v9�ť���mY�#U�D�uJ|�����#MR��(���4%_B�>��L����/knnd�&�^d8}���yud8r5��ud	�n�dl2�n���<ր� @c`�t#�÷L
�cEZz��EER�.����J��@���SW|$td.9ҺD�����\v!j��#�ne� @m !&��|\o�A�pp�p�J��D�\ᨹ�P��
����x��z*� Ub�� �y�*�&�A]����xE=�%D���TC7��xyX��Y�jЖ��=�bI�M�=�5���C.EL���u{�O�>sa�����Z8��[,�/�S��)*0�T�4O׾���˯�٣d�^�*R�ڦ͓�$}kd��bisEH�S�2;��1��bk9�V4��m;0HF[�g7)� +XZ�HD���ިO�ɘb�="sK �x�^��
6TDdu��%��ͪ~�Z��P=7V�Ąf:��e���F�6O�X��m�A��b�����DZ8J�#z�:����s��|�hs,Ǹg/SHG�!����O����G�y�\�Z�9Fc����ir�L�HG��9��_U�)k��d�fȐw����n��]��j��L���OY�P)�$��㗈�ȴ��D��[�5��V�Y��%�!CCb���m�m�R��Zt7�ih@�lHG���x@h�i��-PQU�~��E��%��̎A�EF��� �$,N[`��,]N�1U�&<�i m?�xMkoq�[.���&�?Y6b��aS�r�O^�d�����p尳��H��WL��὜ebڃc�`+��>�Ѿw�2!S��6��� ���wOlHG �B&zz�k�ؾ�UL��:�Y�ci�4���B%I��͐��0�r۷�,�y�5c�#��ddS��@��T�l�vvӣ�}�3��m��af&���B ���AD��#t$b�j�0�=S]���7)2���A>E}d�"�� �5�&��dx���<����o�0^	�T��ܑN$��@