BZh91AY&SY7ʊ �߀Py��g������`	{q�$  �Κ�Q[5
��&"zj0��5����mFG�I�h4�*T`       ���a2dɑ��4�# C �P��������@ �h`LM&L�LM2100��&=O�=��MC�zF�z��d4�h����TI�)�-^rZ�#��*z*��	H~����` {؅�7p��F���.����嫚\�*�!s1Us333332��ffffffff.�t���.�= ���{x�S]�`дJ�лv�Vw�P�K؇�� D`�ԝ��an+u �Z�n/z6ٞ���Uuq���	^^�p�D��������1/�qaR\�ܙ*�Y1�4��ek��'���o� �Kj�)�H�9֭\&|�}��kU�x�hdJ���E�fFJ���%�ʄ��$�cEUD��L�0������2ggw������A���jku��}9[�&���Y�6/�fՅ�uf���5�yn�P$Ñ���r�yN5�Wv�x�%^<�a�s�rĞƉ�G�D�R���T�d�� �� �(�X�qݛ�3L�Ћ9�BqL]���rб�)-
E��K�
H��+�^i�0�p�!��k�#!��:�"rxPӶ�i>��L
'�Z��tSnl�3lu�㈒���tGB1�$�SiqTuw.	b�.�h�,o���)���� f��fr	(OC\q�1�S�R�H����jR�"��% �C/楶^���ˉp�	 ��L�V�Ir�j4��CB#�bY���Ƴ�M/��#J-�}*�L�"/Z���	M�)���:뀕�uqKz �Ö&ynǐ�U�mۑ�9��N��E�}� ,+����$�C���T�D��{��(�ӺP��I�f*)[̣��������rڐ���2�������V����w1]�s��I	T���P��xYi݁V_����9�U��q��#�z���(�2/�!r�*�
�t�ȼ�g{�m��c�4�=�0�F�9��ހ�J6 q��!��C��W� -s���sӜ�`yOiDQ^�UA�#Bx�����0��+T�^�P7n�ۺ>��µMP��;�c���F��T���eR���1�T�J��,X�w�ܳ�j�TH�6��䘄�j�$�(KM��V�TCt=�m�x���͆�93�x:�Y$S�+w�Ow��4�
�v��n�Q>0�_:iS���
-����#���]j���o(�O'�P���/+�R��F
��������oT/W\Õy[�2"A�g�y�٫̲�Aښ	�h��|�Yn^���<h	]ʫ�Pz��6�0�\�G���w�y�}�i��F�E-���y>��?�-ms!JUZ��JïlM��$�#�rK�λPŁ6��@X
Cq)���E`�i�01�mn��eg�߸f���3��y�Y2������1*b�@�dx�cK�L��B���Yƞy<gJ����ʌAj0�T��_Iq�4�/��f�!��m��i�I�~��	Ͳ[�#F�e�����/z�W��kY���s I�����X7��Z����[v[��2d�JG 	~���&�e�d��"���.zM�x���.sK�J�b0Ö4���!{F�����Y�vF-S
�T��B�������&g�W85ĭ(�(M�w�j�2v�C�VP���x���\�:.�aww��+�� ~y��n;��[��g�ȁ�v��w����9|d��m��0.��(�2fh�������k��]nR`��L>0���+��s�Q@�EA��P	J�����.8��A���P �pӠ�xl,`rP��	$�Z��D�=?�_��^�8ʌ�	��d�+)�ǰX��4EP3����dy���Se���1����@4��5Y�rE8P�7ʊ