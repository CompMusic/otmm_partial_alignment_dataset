BZh91AY&SYẠ �߀Py��g������`��_u �0n{m�8�+vu	" &�"=L
2z�)�z�� �4�A��QOMF�F�     sbh0�2d��`�i���!�I��jh��44d   ��P'�� h2 @@� H��&�*c��z�?T 	���SCN��ݬ(��)P(Hq�
άd�&�8A ~�H��N���I$��y/E � *�e<�����z^6_O��ǫ�m��ݽ���mUUe�UL��e��6ffcj^��՚G�0m���V�+OO=Hk���q.%�����f��5b�A��W��D��X�����v?�fk�8�,��++b6QUs)��ic D9��4�4���%�t�6�Vo(|��A���Gw���^F.A�֚�`o�qb$4('�Z�
�J������ٖ��A{�6Z�s I�1����/�Л��d��-c���� ���cK���L�{�܂Z�PT�u@`ň�]J���˖qQ�������d8��PLx7��ZFf[� J��ў�^�7�"�qx�""a�;!j-�٧41�d̲tr�� =�J��H�4mHmY�zQ���2t�n$����17�9�����J�� MQ,�)Q�Lp�_!.@��sm鹤����.�9���O��Kr�0����QJ��X��r,P��L�c]���nK	ɤdm��̡X%���.9)V�Ïf�O% S��"_'E����ZXv��WW`���̝�5Eᬽ!��b[1��p�A��<6�p�0�[ �0��h�R�.e갽1�5:�N�^$�L�w"�`J�Ѽ6u���r2Q!�7A`�9<X:���0df;�����H��}�)����O�lGI<��ȗ��
���S�ѓ�[���a�[�lP.�S7�g���E�'TJ=0hSGfd~��� ��#������Or �`��ؖ9�FWS
�ѪШX7�,��Un�A����i��=3��Tm���&���������fW\B�\-7�������>_����4ƣ^Z�)��0��!��(��U��	���rv��̯.�0$�ۚ��j8�%�P���,�JYuHŊ*�WFTm�2S��b�S��N�\�S95c�!bBf�a��)AQ���vn�ͦ���D�n}F��1;=P���KK�O.:v]�i�7�Ww�c�Kg�|������̥�l%y"q�{��hߜ�^钽�أ�f1�h�k,�̈́����;�-�-�H���3Zo���J�"�h��|2@�ٕ����@�]�l�{��?z�'O(9��|�����ћYC<L\�Æ#Ry��b�����Әl�[�W�P��ET���Ȩ���X8*�$U��b
 �n���0�U�C��W�v��K�H!1G�h����Z��"���	��y��!ܠ\u
��.B?�gʻo��%M�H-q�ӡ�%�R7(GI3_�:Ⱥ8�`۰�H`UA�^U�f5����J�X�a[O��ݵ��>�~~��ٞ��	%2���&���i� ��a�+Aq��	gH.]#J��RSՑ9�@�4�P+&�Ġ��P{�ۂ"����(��2��g�e�����s�(d0�&�Ӗ�^�-8K��X�N�w�g+C�{�V�����?Ӝ~@ߴ�P�5_�ҠBX�ĺ�BKr�]Ao(-	��v���Q���i�X�����b���9���tή�~�h�hсb��R�����ģ�D��Z���n%�F��[�t�d�%��H�O�������MGI Y%�,�D	gЮ[�����T�!*�����ۛ�k���j}�H�C�"���)�� h