BZh91AY&SY�kŽ 9_�Py��g������`	_y�j�  �}����  )'����ѡ� �  ��!D��15 h �0&&�	�&L�&	������*OҞS�h���ji�4���@"��54�6�'���F�  h�AB&O$��2L�CA�@22eTS	=��B��^+������)�`z�$@EB��/P�N$	4$��Kވ(mEP'�� ��t���'t�x��ݬ�̬���l����[�8���Ƶ�W�K.	2íG6����PyS\�i� �-�8vU��0@8�^�!uX*ql�n�
m���$� �NQ�gt�,����P:�����`���ʾw�΍����@8@���Qw\�ڗ��n�H��*�vXV���3�Y�"$
�J� ��#��p�;:�
L��C�,����/���wl��!���~�bA���&z�옘��6C9k�� fމ�� I���ѯ.��⻇]�i !�aݬ�b��3)Y#+B��)(7��]0�*j�WLh�hFچt����zK� M�!@�
#	-)�:���
l��Hō���iGL'v��6�vC����%4 ,��7{����w���p8wh٘�E#]X!	��KE��]9[0�EXfuTB�5y�������P�� h�ҧ�6��y�֢T�R�����h�I�Wk����~�ǆ��Ξ��l]�x�ȉ��f&U6�<@�������LL�_4t��pt2;z�b/���d>�L�]��u���h$ӱ�����.F�+s�z��;�NmD���D�U�0��y��m\�qzwe��[��5��/��Za�lL�Đ�TҀ���Q�9,,�.� A���_B2P��y�Մ��U��i=HLl��3uKr�Ҳ�8��6�{S�#~�
Y���E�KR�@P��5M��֖�b�i�8��yG��(�*���Bw���풘	?��[�̙HA�da��.��;�5C�4)�3
�̲�є�lE o��E\�I�*[,\Uj�ޡL�.���j�U���.��r�7wIꭗQ�7`xY{0:	�`�}d�bi>�or��M0⫖k��#���ֳ�ܴ<�X<�=�C��j����AX:.֞��ݾ~8`�9�JbJJ�j��whY&����ӷ�F\��,�(F���B�!�$|@.j�U0��+US�A21M&�J���S`1$I�`2;"%�X�r{���K#n�8F����S#�V ��d
�`I� �O� }��]�5b�AB3�P����]�D��)�ܽk��&��)��iY�_ec)%�������|8�FT7DPX,��DQAA'��@%�n ��遛�/������'���%
W"!��&��v��߬B��97��܌1�^A�`��޻�l���9`Qk�ɥ�0�ީS��ÿ}�	 ��J��E�毊�
|������Qj:<��U4 p3���..��������u�G�a�n� ����H#a�h���>�̧�v8���:G�]�N �y�y�ʌ'H���1 o���v"'��k !]��v��TL���abL��^�(J�H�+��J���(�\.�ԉ&d`V!t����M	Dn�?i)�[wTM��X8�N%�H&���Bx7��D�<���G�Y�����:n�`İ���ǔdiO>���J�h�wA [��u2�c�4�����>�x����p�c�>`n#�c�7�JfrD�/�BmK��*0����2Et�}r�$.�z������3%/8Zفph�m�.�K͈jC;VI&��w]F�A�f^�=��+�y.P"Ij_%��Y�|o ��&�Q>�����Qژ@.�������M�j ��n��SLB��������A� ��7 ]��ߏ�.�p�!8׋z