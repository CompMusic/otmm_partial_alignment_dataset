BZh91AY&SY|�($ �߀Py���������`?{qk�� ��b
H��&M�����(=OHd2CC#i����h      `�1 �&	�!��L����SH�2 �i�!�    � �`�2��E�F�S��&���F�Ѩ Pjz�4ʢt���!a ����'��-?i����^�>v }�BAr1
\�B��M��m��l~=Z�J[k���wsv�����wwwu�"s@a!H�o��*<�!�6��aJ�	��#Wl����4��,�F�:Z�d��v��7R���?�vO��C6?1�\����--b���T���Zb8��n�l��,��˚��&&��vk�@�����M&~��2-U�ob���!i��*��_y�tSB��
X�bܔR�&��������E!��<\3��i���kf�>����p���Y��YLP��^���[��%�L�լ嵒02!P"P�G����w0{�k���.�aF��!�l:sw]��@W��x���J���� ��v9��tC��	�v�t-�5:��JB�U�4�!�C�8��⬡��I������zXr�A8F�.E�=����NŴ�b젣�WS7;d*cVaY�Hǃ Y�|
�&d\9n�U��#g6ԙXA'*�`��-$i	Ey��n{G�J(ӵ��1�������
2��@*	��'���^���
�Q{�X�0��#�k�_O�h�C���$�3²�b�����S���a�鬯�P�-z:o���!ē4��@v�r���b�P8����Ȉa����؊Q�0� H�T���tcs�i},�fN�Q㾰�Hp�������d�ې��ё���Q9���"�5`+޸w�p�;4j��E:� L�0�:1�v��Q�t��uE�UTH4'7{�r�o�f�
X+iE)3JZx�OTZ�i��II�?X����3)K,���+F�-i��7J�VD�`l�YHЈ�lT�mbֺVhoS	��k�E�MDEV��M4g/;l0!�8%�:L� f&ʧ�k9����'++�]f�B�<p��Rx��h�ޠ�l��/}G���U*p�z�4�O�c�Kƨ�7h�G7�SM�u��$s&�R޹T�i�G�Gɒ|��}����:=$��L�!WI��~�6��j�% �'������6�}`��{���y0�snۻ�����Ғ�|P���ľ���I����:֯���Gg:���$9{g���E]���7���xq@�) ��ib���d�\ၐX�Q8Ax+^�d�'�q}rȦ�& �I�f�1��^�L;{I��@�7Wij��@�
]�.Ja��~����w�%��E���ڍQ໊��Q�H$���"���_����H��<N2%fܡ�ظʱ�mK20��$��O}��8]<uU�����$�<��2r�E>���N����H��t�觸�p�Bd��W��S+�""L�L�,P� .�}�Y�9A*��(F|�b(L� D
��a,��p�;௦�w���X:bsE ��W�A�����*�N�KD	�<8p�|n�8�܃�Z��8h#�]��������"�n�L8���NAdR����0ߖc�ߓ�F�9��wИD0�BL��A�	����ˈ�P[�4�g��U8���ؤ�A;N��BD����80��F�B�@˯���|5r2�RKR�P,�����u#O�5����c���4�[�؊u�5Q5��7k��^h���2e�~!���LD�8�U�ܑN$!J	 