BZh91AY&SY�˚7 +_�Px��g������`�,y�g wa����p�D�aƤ�%4ښ3Q�F�@i�JjOSOS@h   �4�ɓF�� �0F`��T��m����=@�  4=@4�ɓF�� �0F`%4&E6Sb��hi�yF�4�S���"�^_0"XTM!� P��e?Z�"F5��q���� ����$�.pI�V���r����s�S��8�%������1�3231mr��ƀ2��/�Y�z��k9��9�!�b�����3tV��n�oaΎ�:��ÖY`�T��)I�qkQ��5��E��?��f��	�\x�}�r�%�t��:P�9\��8��Iu�*�����h����y��T��ʥ�m�~�.\iT�^	�n�\9��TӺ$R%y�4V���&et��[Ԉ�0���vW�)d�k��.�y=^��i�j\�H�p���7z*VkF���[�k��m�Zv�S�궤�@�7+cE�)l�[��5kqtWĐ�%p##9�^���y�/|T�%��!���=P,�P���� p�Z��[M��`����CF�)%�q��,�%Z|T(�tfAcc!n�8ɵ�`�XP�&��A�G")M��U@�E!���B �#7:46tE6�xcr�������Q��ꂄzV0C���Ra҃���#Y}���(�3�la�����9�0�o����$ZX�w}��}pFS�F���B�`y�my�}��������}��g�Qo�C�*��l��4+E���{�=uSΉ%Wc�D^�Vژ�J�p�45�S�j�����R�(�,�>��鼚1��m��D���R0#H���(��Ƌ�%\�#6�]+	@�5b����������z<�HZ(�Qo,,0�i3�: ۬B>R�pE#,T[PeAa���"��0<!S}�z�cf^��� ����Ey*�	TS���ה�4u�jf>��2�E,��v\;��+ԍ�1|1�G�&a�`�	l�B��UhJj�̻�r\��Gd,UK���`vH+X�����M8k)*K��D�%'��tףX�.��,�܆df$�nupu�n�����ʸh�������}��Ўv���Ck��۬�j��j5�U.|?=��!�E3={���{��B
�!w(߲�pe>j�d�>x��
:�w��	�����;��3��&���2%į�R#���Hp8�zw������ß&�;3�HB��y��R������������Aʨ����OL��'�����I�(���	�u;�t~5��v�-iZhD��I�I!�D��n;��#-�V��[�� �8��"-��J���*�i�0�߭��E��[�����Hk��pb��1D�JM���ڵ�7���iL8HO�X��(Z�$a�-[Ue�A����G���ѕ���6,#y1a�@c'V�'��\�B�9HL5�9�t�|+�MUU{-ׅ|yy�@�	'���ۂ���&)Cܓ�3D��YJ�J^H(��:��qZ�}�V��a�����:�Kܱ��bQUPB@C�M��K��t3a�-�zb����4���T�~�� �]ɽ�:�%�yz�Z����h-��(����]T�z>�r{Cg]���F݇Q�Т� �NS�z/B!!Pu�!����C���tQ��qT�9�t�~=�g���nQ`�m���>0��3��B�Jx��qB�*�*٤��t��eG����^�Oa�ll��ݍ�ZuV��T��OG4(��������܈��10��4
;.M���6��t-璳�pЍ~��'l�+�Vo�X����H�
9sF�