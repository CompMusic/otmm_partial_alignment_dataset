BZh91AY&SY�j�g m߀Py���������`	�z�q��� h�t�\�vݺ�`�!4hF"b5CF���@4�4 �JM����M4��Cs F	�0M`�L$҉�!CCC��� �� d� �$M��4Қ?T��zC� 4�4��MSɊ7�h��&��A�hJ�j�$h��!��� T �_�a�̤Py�$ex!��E�wA;$!\��ə���<x�_����Ue�wv�7�w�Wd���f]��Ue���Ћ�Q�M���p����X�^��`����$�2�q%��Ţ%aó�=�I�r���.	$a!�d;���ӵ�=.�˄�T�D/,b9�q�=�"c��4'1
L�fw̠L��x4i!U+� �z$n��{�T�kE��\I��R�Q��O(�s�b|$ؓ�B�98��TDDg��/�e=^�`*�	G��a�����Zg���d��/�U@��{]��Kk�XaB�E��Eϩ�H��Q�L[��մ�Wj��Ԣ�Ye�+f�$ƕb�oyZ���Ȉ��X���id�g�� �LE7`�t�qHG]{�a��������(4I*>�(���B^猪��w~]�PPQ�
�f����YX�;&:�=ANHi�f]��VJ�bauw�a�>��OD�A�������D���g�!%��V&�a�� ��V"�B�!0e���������8�����v�2I���U����(�K��^	ǚ%�2����Í��Z�pm ��h��P��<�x� ��"bU�y��y?���c�F
��d��	�,Zǈ�v+J�W"a���+t���]�2sG@���3��::���F�#��E�<��KT����n�aںWUA�2���kyz7�]�n;Xx}Ħ�p�W��?O����߀��4H�wQ��9%V�[����5�`�v�v$m�Ƌ���7E��lp^�gFҷ�N�� �l�:)��7^bJ�hm�JG�~�%�""�#�ԙ�s���i����*O��X�]�c�T��x�* p�x�1aX]nr�nf�]�Q 5�N�Vƨs������\E� Y
����obc�TS��su��;͹y�u׶17� |ǲ�(�yU�*�$�ܝ�a!K<���uR���Ee�>ٵ��T�(ƴmij(�k݊�LUe�Fj�d4ٌ%��M�R+dUXk#He�(�#*X��L̀�T6��G8��..LhQTWf�Ț�dw����ن�RM��jvz�ANr��ٻ��Z�2�����Q�C�Wu��G��`ϛ�@"6�<��7��]E[�=Q;:�*�X��f��6i�Y��'�� >�^�d��4!�=�'@�ʭ�l��;D@w1���=I����r]*���	�u�^3c�a�6m~
�^�r�⹗V�{u��1jOr(�[�K��QʆU �y�C��/Lb��^��w1��Md�U�v��D��ӥ��2r�I!@�AH�1�3r�*�2���2t!�Aۨi��3��	a���G���Z�
�TRY�	��/ras:��BVhs�	j��g�Z�-�&h�ۻ)D���~o��I{�:-�$aU��2���0�d�(xS���gXW�
bt��z�#g�n=�	���Ć"�/0ԏ&g�o�4K�b�$����I0����鴆5��q��[��"�̢�P+1}���$&�r�-Q%Nd��a��� r+�����UrP�8!�Y�[�$9�I��@$c��(�*C#Kh��H��	�rq�,��)�E��Q�uj�\PU�P%��S@�^̶B���� `���]&A�ggG<��f8��<H�$]�d5n6�1h��ȉ�A ]��*�j:<5_hY����9��P�d4�]��x����3��k&��>3ʓ�q!��aJekf͔Z_`�R0.)��;3�ۖ�*��"1�0�]���amX��KXI'%n@$'�'�\Ю���g$����AuZ��F�W��)f�<fUo&�UY��L�
�DY�R�-�����q��z��-��.����H�
W�