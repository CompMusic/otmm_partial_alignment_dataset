BZh91AY&SYKc� ߀Px��g������`�1�v���t<˻���)P�)�=&��hh(�=C�m##�4C��i�JP��Pd M@1Zz��d��Pd  �� ��!���4��   4�ɓF�� �0F`" )䧀�'�eO
h  ��Q�����"@JH�I\�(I?_���2�M��P�0����� �͖�	J�S��xO�׸̽��������ݙ����U3�U���
C;~��TwÇ��;�N��[,V�)e���S�����@�9��SJ	!I���������@Z�{ �P��͔�+����"hfeyD�Rf`c��*%P�(S�p�������ғm ��Q H�ao�1Z���UKҿt�iV�Z���d��fo����D�E�ym3Z ��c��~�`����$��,M3ix��f��AkHcM�3L�bT0��"��Pݴ��AK��C��X�G'�5WR9/`�)
��J��jރ�6<�%�{.�A#MJ1�JB�M�������̆Yi��-���.�!�� .�T��QN)�f*�D�J�j��b$K̛(iPӑ����VJ!Y��rX(6�C�Z`5��]Lcm����	��$c�eE*f�PbE�����&
9��^>�Su�9�����qhq�w-/�E$�J���������'�6�yJ<(��.�A�UONѦ�ъ��]��\,ܶUJ��\8&�J0XLI�ɇk�aeX�mU���X�7C2�c8���|ָOF�q�u�劝Q۾_������k�B�Ej]D�rg�p�4|�t�t!�7��
Z�i-3�i��bGI����"��Ts�����Q�J(X��g��qZ�VVY�� �e�M����!p h��s!�.^$V|�+R DD�;�(ہ~a`�CAq��Jm2
E 07#W�!���N�қeeN�P���R^��J�������-NV��T����i���k�W�Yc]7���@�7\k���!�FV�|����;�Y�����/KF�{݈u�|]��7K�5�.J0T�Gz���~�/�P�/$���@�z,�G���΁�WE� u#v #%����ۊ���=�:�O�����ĈR�5���ÃGn�!,{1'�'��v��Z�"w�I�.���/d�Je�����6���K bcm�eÁ� ��!P��iױŌ���SH,�b��FFJ�#�H�ДD�
��3ج�E����{�l�����>*ix���Q���]��Ž6X� �"s�H`x�[�DxY�+��TOu
ڱ��������,����0<�fB�C^G�l%tw�i+�k���M��J\Yk�3:y;���;���:�.�����ȩ�x)�PъF�͠F#�4�f��	�����`���l]��H�+�	�6�q $��ä։���Z1`U�g���/B�#2�!�×�������4�Q�ᙘ$C����H;p�q��r��Q]8�|��(���%w��c-9���>�2�0��z`�n@�:X�E���%d���L�5&��&Z���v|cb*�u8��l�lS�$�~V���o�DM��Z�����$0��,l������lJ1�q��jF�˃@�ϼc>`�7*Y`���|����n�n@�;w@j��h��*���5���3�y̅�j�8X*v��ܑN$��5�