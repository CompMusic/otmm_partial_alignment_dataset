BZh91AY&SY��@ �߀Py���g������`�-��΀"��VJ��@B14�F�i���1CF� �@�4��i��LM��ah�0`��`ѐ��&��MI4 Q��Q��h   �0`��`ѐ��&��$�4�4�=&����z��@ dѓ�l�<"-  ��E[ J��C�V� �"�u�e�xۊ� ��|��A'8(e�Y��W��hӪ�{*��hs,Ԇ"2��w�O��Iy$�b!�Z�Xii��W����K�Vv������]�G��L�>��!u�Ѷna��H��CA �K�;MU�-މ��  坵]E�pv{��20��O����;Z�4��h�H���C�2D���=���|
1�$�Ǔ����.�<=5Ä��@^{2圼�OC(��FRr�
c8�,�RYB�8�ĆYQ�Q�A���jq��esՆ��7b����bꃲ��0Қ[��،�垰�`��8m��1���p��-����(�p�N���$��(�8 �M�m4e]`�)�k�"�Y��K/�&*B�hbWhp��Wp��Zi,�6Ȝ�/��q�g�#k��L(9q���a1s��6�h��j�[��E��Adp�%��H`4�W�5T��`������/
 EY �m�⅐6ק�t]�R�旚�N�am��W!a��T��BCl*fKȖ"w��L���J"��*�HЛo�;Тeߟ�cfָaz�����]kT�7K��UI��	cW$��,F�`�b�˖�X,�C�T���)V1&�gP��bA�2ɝ�p%�L.!�8��eAd���Ek�Z���i{�%]\WWʠV���\��&?�w49���$�RIo������J�	:���]@��)���_��R���Л�]к�e�}�l��@7���ͻ��s@P]�wg^i�m��t�[ Y{���P�ɭyd?��g`���"޺v�HW�ɚ������p¡F��-?\	j��)��3c{�g�$�(΅)$,��ZnN���ܻc��[6`)2A�H�ƅ�,�!sT F_9Z!�/~�c�&A�;����d\(�HB�%[�nr���s�i��8O�y!�j(2�a��iQ��
�,�<���޾����E4X -�T�O=/������[ːO6��l*Hɝ����%�_��D��[�6��֢�1�f�ቁ&�?,@�o��4���Փ*����7:b X��Q��0:��*�p��Zrj>��.�&jo)|�A@��a+0�g��Qcl7aAwū�a.�(���� /�Mľ�ɻhja�/ۄɻ1hu�&H^M��p�M�?z�n&��ih �>{9�{�[8e�lA�`s�����O�7r�{�Do��@��@�A��8���bun%��N=ׂ�@/�j�I�	0i�8g'�����a���*2�j���m.6pck�����lң�+7��^�+��7��D+����)d��.~: D$��g�CY�9�`/��R� ��TC�G�7�́v�8���A�p�Oi��PӠ�}�V��[��,@��EO�]��BC8! 