BZh91AY&SY��\w �߀Py���g������`z�c������fj@H�&AS�h�J2b1S'�2�&��4 "Rji��`M1IS򡡦ɀ� �0  #	5�� �     ��b�LFCC �#	��d$��2F��=C��@h=M4ڗ�@��-����� .A�4�!װ�~��S,�� ,$H|�_��!TbK��;F�JȄU�Yͻ�v��!�������k.�����������n�h����Q_T�g@n[�n�em�v1f-�Z&4�M(D���I�E�D��RY����D����V5絍����Z�qqqQ���e+�.ge����5�Ħ�}�JVJl�A)&4C��&�9�E�ւ����
B��u"��`��KwG�F�luܦwCI�%<�`F2ܑH�Z°�s�P��",UV��ӈsCoG���3,�ߢaG��D�*8���9�
�N#�"�A	X33++���pP��3MZ(_Q��r�s�����E�8��1�PCWV0����mT�JsK�Xׄ&�lp�M�*Ҷ�)&#C7��%��cÕK[�7+sy3��tsx�^�6�WҊ?�f�]����&��O�p���Gb6-��ɢ�*.9� �a^�D��5E������>�_���սA�Ԉ!�YC$��F�P�n�.Nj1)xƮ�-i\�B�"�T:8Z8G���zP��PRF�p���Y��(xD+��N����Z�zy}���ք�`ʕ\V�<�7A�;qZF��L����)�Y(�pp͍��6bl�ި��0��5RbٙM=�K��i�K��V�53�!r���2��Ѯfh^�g�!l��)omzX �>�l �D����&9����Bp�g1�
7 9;M��y�!;>�*�8p�����хEu4@�H�TC�Xi�J�էc��u�ExꪬH4'K'd;ШjpJ�?묆P�o#��]q�(t�ұt�]�mf���3@`T����%�e6X�uI)6i��L�Tt2��`D�L�%���F����5�J'�՝]0L���Yћ�B ,���l{��{��������9~��}���gmg��gj��0j�f
�����?������A���Q��걖4��Q�^	">!-z8�.�= ;��BEQ�l<�p}A���Qk5f�kk�q��$i�mպp8��j����E��q`D���r�ߛc.DZ��#2^K��m4)8�Xn)��[9�V������K�Fӳ�8�J��2��/�v7��,3��E�
1"�ƆI���=H&���qk-js���RE��dʏ��β�)�F� ����*�X�ߨ�r�?VN`�Ppj�@`��*G1E:�r]�JP?��q��� Б#a�A��8Y�鍛���Fa�|���I4�;Yo�>\��U+����lC�{ܸJcJ-I�2��mІ��C���k^��ѱfh������]�5�9DC����G��h-E�X��I�!"�(����|��ei	r�Z�S�J��H:��c� ��#�!M
�*M6nL��dRh�I2ra��(�'6T��ԓ��A#�.��<xƀRb�}��v���a�qH���3v���`D�����p�$d� �ig��F�H����e�o.�����/u��Pl�0߼����\�η�FMYZ,n�IN��$n	(b�h�$X4�с��Yd7ϯ8@�gp�,	�7�C}���)+`�PFM�@�2�y��#�>�i2Z�# H�B�+M�P��h�$z�B9R�emf�eYe���G0�u�"l: "Y�_�]��BB��q�