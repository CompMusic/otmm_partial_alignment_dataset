BZh91AY&SY-�� �߀Px��g������`	?}����� �Uou�wu�<$�M4&�#�=OQ���=A�M� H� h    �4�ɓF�� �0F`��F��'���4  �  "J!��i����ɑ�� �M4E�5@h@ 4  R�%�T���(J{��alY! V5�Ɋ�U@�D���(�f@�n8U�=k�p��{i˝�F��233332��fffVb�f6ffd����̜�;��B��3��i��ׂ��\WF1 ��a�1b�3�`���sla� �fJ���UWLLK��2츹eT%�yUwъ	_���(|��Hv;!�6'��vW�vWa�k�G��F�Y)awq��<IV�	Z6{�ex_��Z��+}|�H�:/����̖j��^xk�)ivI$ѡmW�;Ī�$�rl{�4�U[���o��=���^3מmzhq�m�,G˙1H��UW+%���x�L�K�:&�{�Bզa�7>��+E�X�O{p=Z��*e,f�j��Z:�ne�	��E� �2�<�1j,�JR��Ʉ]i�q�t1F$�
��mGAl���R��H<.PP ��o6w%g)%� �i0�rfaK��9ƈ�l2R��K�
&�wTr�㹬I���Y:%r�� �|���CB�@h'��ӳ%\mpɲ���l1J��N*9@�U��Aj]��NT�4�fU7�6��r.n8ts%��5D���R�I6C,GGƌ����迂u�s��W��a��;�0 ��zB�FM�T%�`q�U�nh��D���$����`�n��Z816�{RՆ쵈]��\�h��Qx��T��6K��N�G[�5�J	;��T�,\�����IT# n��Y1i��P��9��'�DDxqC��c
C�C�?�B�w�2��ܮ��
�:���5��%� cTA�V�J���a/F|�H�(�������C��ؐ���mJ^����0]�p��/.��o�y��Tp�ڇ�_��(�+�UE 'o_xyH�(�<�7oy[�UT͎�}�۵TV���E^RU-R��KhZQ�B�V�Za�AQGd��R(��L�Ɋ��]�EԘ����m"�����l���3+.˖%y�w�
�ͣB5�^� 1V���&��Y�o~XyO|>�_��C�*ih��(X�<C��Y���嶪�kI��~�����a��黥�W�O%�N+ܯ @���`2��������� ���B,��)�eӺsi�x�U��@K�į�UWVǴ��d�@c�r�]Ip�Xu�ſ�2`�Q�"��6�6������ s�$۲��a����ΕS�I+OVM7�k�L�=�|��~lffKxB2$`B,"����E�QJ1��h<��zL�AM3M�J����f�ZU_1$&Q��҉���%X�<WD�#��b�P���!@Ej��d���@����׋>�	 
0�@*��rG��rث!��%El4ǁ��������q35�I	ܘ��W�o,��mb�I%xf� �b�w�P7�yz��ެ�nE�s��@��Z���<�D��/0����,U}�WL�n�t ��v",(  ]s}S"��bl��	I�2�A"Jε+����@�+*����Nt��Y�j`��م��J�^� f5�y2#5o&�V��J�0\.�~��h:sâ%��*m�����y��X�=�#zp ��A� ��
^Up�*�\��t��]���M0,sa�F֕2�<~2q�X>^g�������i��E��Ib�cs�uR�*j�o�I)6��կ��TQ�ͥB��v�U���qs$�rP��	$�^��-�a����M��Ţ9���$��J�^T 4� ܜ8�d|M�Tb�2�g�c���GFHSx�,o�]��B@����