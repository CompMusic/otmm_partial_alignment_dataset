BZh91AY&SY��'% �߀Px��g������`�{q�{��0  �U��։H�#AOC@	���i��d�CM h�A��R@       ����=F��4 �   �P�C@ 4�   �4�ɓF�� �0F`(��*~�A�=S6%SM� =OH\��O��Q.TRȡ�@(<���2�T�$eC���  n�!K�0�$�2��mmi5kٶ��uu�q��2�����wf���/1r��@4����.�= ���\nF�MLC-;�u���wz�z!i�bC>��](���ᰖP�)��"`�M�$}ͦ=�M��ŵS ����\�m�y�q�����\WFD�\����aKZ��Y��x$��<,c �+aU	�s/��e�SZoԬ�z��h�O��H���sb�%�i "8�̡�Q5�� ��$�r�<!��ҹ�:i�����)����2*BM�t!��Hf�J�m��u	*� DUf�����0�ZXX�e�V^A9LTm`��f
�
����r�.@wmh�<��5�I��( YN�8UODz(��:ʨ:]�#M��+ �V�8�ԫE�!K⣐5�riX�ņ6��!��-2�؅�V��uΤ0$I7�Ä��`C���V������"{Qӗ%��{��k�Z3��⼔��6�'��%A�7\�E,ь�:�Pܤ��7��6�1�'P��E��"�V�,��nJ`� �iNPfE��q$K&�u�+,�P4r�@u��H��֦T��u=����x+n�e��2��"+��s#���S�;,���/�)���l8]�֡��^�qLP[
ܗf1��w�6��

R*�᠆�b����T8�aD�]�İ����礦�rU������4���MP뚭�z3f�8�+2b+�TN��NFP����aHk,P�}YL���@M��bT��3*�T9�?�r��w�ZԝQ�~���X���0;���(9-�da�#iU�#G���Mv��s�+$	��hfSl��,5F�96���"��^��+"�e/�� �A'�$�H H�?<��7��8�gT	1\:���y��P;ma���cmi���	rȤGvGY��k:�*�G%R��ճE�"�,Z[EU�k*+�L5V��**�͢����"Z�6�y�r_3�y�t좲C1S)���]��^��]^�wpT8u����'�i��x�Pl��^��vO�橰j�����:�X�=w���Y� ��?z�0�T�˫���K��A�/B�G>��E ���-���7�px���(�gM= K>��1�xl����p*�+�5?�a�J�T��C�e_=,T�J�C����Iε��e�d(Hzi�jR+��)>��X!U�z�O�Y�Uڐ�PE���hdX�5J�a2v l:�n�ڙ��� ْi�̸ȋx�)W�,�umc�n��� n	�.�Cqb�f�X�آ#��X�s�-آ�pd	Cr��nF���d̢7��B9��"+�+Hˡ�sj$eZh5��6<a��l'�t�� ��� I���Sg�@n6���e���ץZ��6��I$�i.�k�G_��,����d������E�\�)���2���sـu�^_S~4*��s����w�-��'��d�Í[��aw��s/�;�%�,.�'_,A6���u ��yzN���âaۑr�x�䇁�JM۾n��t�>%M�n�|'�.�X&t�䝠/ ���x��e��lvoC 烢a K�8	Z�P���O��_��ƫ�G��{�t��6a)W�T��;[t�J%y���S����u���n9h&�$�aK�֙m��M?���_��N!�ڻ" /�\� ���H-M�z$O#{}�llB?�5!ƞ5�+�v_���"�(H]y���