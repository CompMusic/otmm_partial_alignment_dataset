BZh91AY&SY�kE�  ߀Px��g������`_{�=�<� 0ܩ�!M$���FL�Ji�$�@ځ�z�OP�OMO�=A��Jj=M4�  � S�P��       j"��� <��  2���12dф�14�&���MMj��Ԛh z ѵ `LI�w�!��@�	�y�����I�B	>��L@	�H�҂�	*��y;�~.ާ���xɯ_ɻ�32�����3+331��FB�&[�����0W���MN���8�8�/Z5WQYN�0T�vvVE6$C7����y��́��!=�^~�A�`��% ��"��*��WP�(8f�3l	*n�$��Fx!,]j��C����y<�i��{"��l�$L��J��YS�˞�Jb�⻝��ը�U��͚�`���:�����-\�����2�����>�d̄/J(�xeo>Dp�e�2��ML���q�H�[4�� �/[��A^xS�JS2�,P,4��Ba�@d�mjy���H@Y
��������J�ܝ�]�<1�0��E�2�mTlQ�v��^W9�r6����ȝ�<XV�5b;%�E�|G��@��)�;�l���TR��Cx�((z���.�����8�(��X��p�I���H�Jd�A0^MF1���P;�R^��ZQ��C�^�H�d�u^���lぇA������Mu)�)=#�f�D+�ËԪ���5K�:R��N8^�N��3��s�*�
���s�0��G�=ɕ��~u��I�de+�-g�
��I&`8$��><􍓦�SڊQ	n�E�N{'6����!��7`^���n�vj3*�v/u��}� �A'�T����=�)�����ka!�����&e�R�*�[L��)lEcb���B�Jp�n�R*�S"�uT�����Z��gGY�t�(�j�/yx�0Hl��#'��e�������w���J�
oOR�a�_<)`ִ(9quq�X��5[�xb�=�)n2f�Q7�d_��`�z5� m= 6�,ΙD�4�a��m�w�	�g�ɜB�p[R��k���d�k��E�1?�/�kڧ�cD�c�_��o��kR��7kb�B5v��JK|����I�2d���QH�A�QPrJ�t+Yi���Cz��p/jI�װ�WL�6*�Ȯ����6e�6J�0hV��8�D=�W�X�����	!���[ fk��jd������N�$'J����He4@�NPU�j��+Ls�K:А��F��5���~�#�u���F�F�H��!���A�wy̹@2j�d�|J����i�[�ؠ�� Z�˴�T�И���xLy�#�
b�W�i����*�����[��a��P5�Ȍ��iv��T�C�?�������~����PRG>�:� �����ޮ�␎�D�L�:�熿U��� ������7n.M�C��&�!�����z���L/���)!�
�"���9m�i�]2h�.E�A�Y�e[��B;�Ր�w\��ԍ���'�5F�4h���u�v�d^	�$A۲T�M���Z�k��&��$Q��?B#�rE8P��kE�