BZh91AY&SY=� 8_�Px��g������`�{q��� �;�q
��FF�M��=)�F�12@4ш4�B� �      9�&L�0�&&��!�0# �I$��<(4mMP  ���C�bdɣ	�bi�L#0���M�S��OM5 i���2���>}J	U/AUY ���%���*����yq���	'!r�S0�Qw
�cy��ݪ�a
vCn�*1�JR�335��fffffkZ������P��.� ��ۈq`��V�,�JE����������ۨ+���r����x�4�CV���hѫ�>y�L{<G����9��]}>�x�M�9�q�8J�33ySik�b�r幘]89�N��O�&�S�wѸH���JB&����X�YTw�;��\f:����+̘�pMƶ*��{�X��{���<�m���|�=}}\�ó_&���ft\¹U�6h���Xnz!:�8`�,��i�Y���<E_bD��]�n��oZ�F�P#R��@��I���_@�'(����Nڕds	,ܰ��;�8q(9M,���I4l�a�i������F�j	Z)�š�6�T5R�-`i]���bC�b���B7Y��XD�Y�<�7[�li��C�g����
��C"�����|�w#0��!d��S�ɠ�*���j]�����+4�n���/�X;����\�,K@d;f�Z݊�d�a%o5���λ�����D(j"��2e�i>� bJ1֣����q��m�v�u�F�.�<5,i	m5 �]��n�8�3-k�5�t Y�!:�*��X��~_'�h�8����N�o9���(�����`���ݏ�F���B�.��za�	�L����]r�턇�^�6|.j�D*��~�]�[xx1�*8���r��)��ST�ޠ��A��9r 4�p�Zq�-y��@�A �㪪!'og|�J�?�]�ћn�#���9O����h����,���h� �i�c�屳p��PXGc�c�P��Jڨ�WCQ�jP���d��݊-�J�h�a�m�x3�z�ޖ���펒L�C1[)<�]���b��g&k��'Ҏ�O��Q�
��7��-�r.�������E�I����f��1�پ��Ҩ�H��w(��䱁���W2_�8��.T!M�:H��c����$��^a��(�$��O����~$�N�w@m�8lײj�f�A'��&P��/����Vb	 �7���>B}wu��{�=w�j�7��p�76�d9u�[�~�rXC���
��*�NE	UT�d�y p5�&�/������K�,�W�yS2��?�L 3O"��v�;�v� 4�]�A����*��^J]���[��`��F��+P�,�)�okv:��B��S}xiQҹ)���xj"hZi5��2��<��XC�KH!L8L6EU�9��fQ�{,����A7sI��BNj.���#F��8���7����b��	���^xDr�:� �L��yǍ��Rր �o�J���(%\�
�R$��"�ZTO�5ųh3`�
���>Vf����`F	���ǿ c��7�<{
�����;�GEaۙlnƠe�oA�ewi��u���p^���'c(�=�� p��:�A`F���[�,f.'@}Τ�!���8��$yfu��(���ut��~]�v�)�r��wn��m�
3����L�$�,��D�Q&��Y��-���KX��9@A'�o=u$_��a����P����mx��^��lDho�!¼�	��_C�βS�AY�F��\?��H�
G���