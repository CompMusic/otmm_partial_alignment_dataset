BZh91AY&SY�U� �߀Px��g������`
{p���`�* t43j#ZU!$I�L���=S���y@� �6P5=I	h  �   �bdɣ	�bi�L#0	5BJ4F�    ��9�&L�0�&&��!�0# �!O*���O�M#����F@��dmM5H�w���@pI ���/za"�$��)�� �B�bpfI��R˕��oQ�v���]uUVf]՛�����Y����̼9�ٗw7mU�wy��#`n���s�H8|�qd��*:�!)멛R�3b.�LMj$�D�<U?;iq��Ά���M��U�T@��f)ŋX���υ��Ԝ��ac]]q�nů"L� P2���li�����a�UE �O��:�r5vG�Z�A�aPS'�������^�X��{�����ŭ����C���	;�`�йM��˜�&�yֱ	������@cl�����<h����1�Lo��B��PT�5NÏ�\6�m]ᘮ*����{t6�w�(���ٝ��L����p�\'�N��&��^��$$��+e��C��+a«>Q�0��vrD�kn�'��4�~;9軂���{��ݒ���hS��l�� �bw��FT�in� +V��.���s�\!��ۉ��3�K�r52��E�R$�m�w9wW�/F��v�%X��0��{��I;qA��x��a��ף�7Muκ���7ah�LE3��v�0�i�ӫ�4���l;h�C�"˗:a�U��Wp�Y8f�n�-&Y]i�Sj��tä�<��5� �Ñ�T�F1L*�g�oCJ�s�x!�O]d�3��s{lE�'p�3���"@��؀�ۘ-���I�w�QV,�7W�������5���ʌ˄�ym��N�2/q&�8A
T��ܔ1��0P7��6.g,L5�nbfy�-Z[��ݨN�4��}u{�D_G�7�]ӕ(J
y�ɷ��jA�CI����~Iz�JH���Жͥ��������Y�U��zP�L�p �2�eZ�D�˱�Øwl�y"���v���`i�մ^�ɳ`�6:n���LO;E�系�����]0�)>ǉ���eho�35L�L	�f2D-���r�����րk�0�v3m}��en����ۼ��Q�-���cA��uCʚ���U���ēA"x��N[CpӾ����j�G9yJ\��3� 낫0!���oDr2Q;�r)�Q��å*�cgk1�5�Z�������UA��|Q0�yzi�X+iE��z�G�� �-F#EX�")U�[��*�J�@ùm4%UtSm4�$�m.�)JD����EX���Ȥ�H��D-5TS���"ٚ�!stb�w�m�*�Ä;ٽ�Ŝ/f쯚�L��YT�d^��ƗB�[_v�~�A���6z3?����:�j���Q�c���=W'����u���ǓM�>*?j��	� �S�(C:{CG[H��2^�Q�}"�x~���(�Ԑ"$;g�o~cvU\�0ؙ�	z��P�lܽ�5���n\tBAN@we�C�x���Fa���+P�� ���zꨊdwcMK��7|!躗�U�M|�UMz䄂Ӟ�jO�Ћ ���\����`�������**�(�Y��@�a2�
v��;���f��.ҟ�M$-�B����;��ҷ�;�,8����mz3�ɎT�P��J[v�������e�*�p� �w�1�Ye�P7�Zg*8�D�ui�~���3]T�ޤX\c�9^�.UǮ�Ԅ��̈́�0�������x��W6[�ڙӻ�T��J�C﷕�&}�#��%�)��;C�ɿa	~��2*�uȨcb|�A�8Dc�$��AK���g�fTK7bֆ�XH�L�M˚N�m1��/jũl`Y �88���bmE;
y�@�`��Ӿ���y3��_��a�__>��9�C2��s"���{>\�N�P�"�\z�߫��4nCHx\�D���I����3��A��[��55�W儎�ֶY7��1�V�cFs$�MN�*�������6�(*d$F܀E'�-�)����CŎe8c]n�Cb(p������T6Q3
��p�Q	�7����/�����A���)���Z8���H�
ʢ3�