BZh91AY&SY�@� w_�Px���g������`�3ãET
l-��z�Vښ�D �4�SOI��j 4� � �5Q�dƐ ��4�2b`b0#L1&L0HI�����2i�4 @��ЍTz�=@�2�CL�i���#)4��54�Si�S'�4 4 i�h0� o�ߥ* ��W EgoaG��$���R4���o�@F�7B��@��,�����O�;���M��K��ffffe՛��z��UYZ�����w� ����8����择�o��W�H�����0֐��"�J���ߎJš�&�|,���sFr��ј��Α�Y^�����ݍ�� �xf�%C��.��{�_W�{`@ ם1��Mx�8�H�v}T�c㪌0�<Y�A��jz竦��(��H$���L�y����BCM1�_o�y��>��ߤ_�S]�<�ʷXuR�❥d���t����b]6��Б`����22���G*`
�C
����D�L%����N��7�tr����Ö7����n�M5gX��$��Oa�Ʒdb�J�3W�5��N�浐� ��搳��,���;��q�K��%kxq-���/i����c��������X��B���* t�Gv#e�A��b��o3U¢�����r�n�a�LO*"�Ȕ�y�o: I$��SR5�t��K`ɩ�Қ�]��ҐX���h���}d/Z���֬kb�jC�×�QaZ�f����MLIN-��"ۍtB�#c���dgu��
�
,��OBMs���׉���v��.}tV��艠���jR_B39I�zܿ�cDRL��o�$qYݎG�u�l{���Vqٗ�o9J��2�5���֭�tD������B��[��K��\mq�S���Ȃ���a�a��a�$��;�Z[z�Y�Uf.!!ʹ�|	�۷�)�a����3��S#"4�B�����Z�x�4'q���ڃ���m*q���s4��
��p���<]23������GQU3��4�����?ڃ���/�EF>����u����=?���(�T��ʭ3��� ��)�"�M���T"l�Li��@d@;J�x\fC���],9I6*��:��\���h7��=���v[aݪI������#�c�w��V,$�x->?)=Y�7���j�ĩ@�6=��ĕ��3��<۩�6F�-��I �RA�lU64�A�1*/��y��Y�1�]{�/'Q�a"U����),��|�2���j��3�RfiA�BG���#4�:�$�֎��dÌ$�G
�dV���G-;V��#p����aZy�-�6�l$��Qiq<�^z�W�[�Y!"�6C�t޿�q�fC��m��e�%�l��I��	�e�&F�E�)JG����v��e"cS1E₦*���=�1�4���B����In�r EXA�v8IhH�����-3d�]v����!�_-E!Xݫe�&|�r)�A��/@'`����V{u/c8�ʃy��\_f�y�/E�,=1�Ӭ�h*`�=�;6�*7��BE������y/��_!L<u,C2h���L�4�z�lR`�,s�L!:�!]�ns�h��=��	��Đ��X����a��n�¸΢�BG9'�0"C�~T �{O;?��٬2W3�!r)����ό�*f�QR�E�:*c�7�oB���[$9)�L�!�����"�(HU�d 