BZh91AY&SY�4� [_�Py��g������`	�z�t�aT teXϸ�7)t	F�b#�5OS�S�Oԍ���G��4?T�M� H� ��    �	���dɓ#	�i�F& �&�#Jl���  �@��6��4�򧩵?Rz�Pi� � SMM�����mM��#@@�d�� AϾ*�(PD�N�������H"�$��$e?k�I���
��]�R +$���������3����g33333332""#3333+1s333+1q���H-���|>�������US��=��9�)LC<��E�4����{�Υh$�FU+\�+(�\�O�t[}p��mv�
�4KQ��i's N�l��q��&��;KuWE��w
Ke$)'c0���N��z�jr�� KRdt�n���wi^�ϗ^����U2�K�-3��8|':.���8�A$���ֹ�>��I4���<x��!7�Em�g�9�K����}�7n���n�Zʪ�/��m��TUeэ]e���ni�NtX��"s�ۋa0�OP,�	�iY�ǱWTa�y�=����z�p���I��uu�ӥ���
q�y����t��z�!H�r�J�a���V�4H]!qz1�t�5�!h2�K��2��:��b��aÌ�ڳ��x���ۓ�R���͊�Ŕ�0xs�M9|��\�Ԇ c����qRtCNՅD*��x�E	@��J`��̧5A��lZ-i`��ч|H����Tb-��4ر�bÔ2�q�#��)�{6X⺖�~>J �U+p�H���q�_�L7/���]�I���&CpaNV��+M�e�W
\�NÐ�@��ք*�n"�'9J�������
�������r�w
S�?�'�X�VL�hlŌQCO0�j�887f��)x״�`��+X5*�KL�
C�W��c�	�&�w�&Z���$�K�`8�ٴ8���$0�5�,Ѐ��p�����-7���j�󜡊�Ö_v���%w���1�{r�rx"sM2�����9����6���˾���x����i0�<�î���Tub��[�$;��[���T����YX�
�3���xlu�ś6VeW8���S�:��K��\��L>#�QT�(��HН�<���>8%L9Y+1��*+ ��c�_3i�R���d��Kh��)
HShRj�AAD�#"��)���uP8B[7��-�T啷IIb[4�i�F�SJ2��T18d�x��|�}i2!���� �BmX�l_*]�����+�����*�ʈ����IG֣�џ�I�U�^frϿ��Z��LZ:h:|c���u��ぶ��(�P$�ɟS�I��,�Q\�����=�q���� �@PKHY�bn���٦��8M���~Vu�/4֟����ː$��v�;q��J�����	�k-���+��^j<�M�4!�Rf5���[�R�����UYb��%����b��+-�z���o��{FQ��"�V
EdX"CLY=&I<��4m2��*l:��ᎃ3^
��e�fb���:Xu9(Mt�8Ԅ��y5�3ÀE8!�FPW���cc��'̄�ӽn]��Pa��⒚N�(��	���-�NH���N�Y9x�<��D�z�׼���A�ʎJ��4b�MqzެǶnŴW���r���<A��K_^c5�6��v$�Hf"d� �Qߘ+�9������x="B�W�s�Fָ�6@�J�IEmy�j�:�E,��u
/�$��xx�a�I�׀�MN|ǫ*�T$�Z�	�NC-aҐ_j7u�{w<�k�:�MEAX)�vq*I=��H$�2(Ix��� �����x����8�I.�A�0�h���|$�D�F��Ex��p!3�S�nxA[�w�'�5���r�W7BF`�P��m6�@kv$
P������q!zQS
6Y��X"XZ@��o.����-����\����(R�Zݵ�R��&� \9�6㙵u=��VK�2Ip^5k���g�01 a�1�e�vh�x�\�^C��CYdWW$V]�P3ф@��0��-R~�LH;����ض���"�(Hy��~�