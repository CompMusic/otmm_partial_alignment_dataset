BZh91AY&SY�?� �_�Px��g������`
���5�d  @w>6sn�sj���50� JoS6P�C��zC �F�*���     �bdɣ	�bi�L#0	4�jh��44�   ��(M�� �4  "�M��4�����������L�d�2]E���6�RH��|��NI��ʇ���Ԅ!����Q�̒7,e�ɶ��y��򳫝k�www2��ff���������ӻ������{����6x�re8p���:E�?����=e>�ѡ"Q���b��ʬ��� �|SFnj.&�<���L���j��-upHZ3U�ug{���N�զ�$�e��G
�S��b��R83�QC<�\cZQ%I�i�m*
����`Y7եI	 J�B؀,��&��i]��j&��u>̕t)Cd���Ƶ���a��C)=�#L�H���L�2Ւ�|���L3z���K���)���Tr�<���,��ђ�p�8z�Q��"���~WlE�� 8� �C�9�I�;��0"
���Ҩ˻�|k; 耓�f��^呩l����*�;*���s	�<.���B����$&<�����\�FW������l."�8^M��.�`�h�S�V��*�
l�(�Q2���	E�x�S1�9n�uI�び��s{3�H�Y��>l�xY(,;$���,A�Ȅ�Y�(³�p�����=��u�V7�y���١�:�DT�^�=6n�\�]>�<�h��e��@�X^[�2r�3�t�1'���T��.�vLGmA<.�K�@q���L'\��<K��e��{�R�y�"�!3�r.�_�l��y(?��34 "�w�y�q D2���96V=w�^sd�#���7B�7)N�J��Ǘ�a��L����*U�<�Pؓ��@�D'V����R�����*h����1Hr�7��7s�3�(���+;�˂�	A?W6xk�ة�j,��t.T%�h��Dp�,�V)��s������[����R�U&�A�u8�ڑQP�f!��m�82���)>���ǜ��8ph?��6��}Nׁ%�@0�G����Q�9�qSc��l8�Cڬz�U�戕ǣ���Ȅ v���|�:8��������v ��gu�^�� E��w�5��5B��0K�q{q�*�+y�L̈́��K�[�/�qN����
{��U��w�!Ė��x����\b;;H�u�7H�Y�)v���R␪��d��|IQS���$�'���|��6��]��ލ�������J ���#EX��h�e�cŰU9K,����h���+�jQ%W�(��*�eTRQEX���IQ TG�4�&�+�$]�YD�0n:Ѭ��TI�Lΐޤ֑\%p�s�I�Q��c��{��i��N��exE�ޟ*YS;G��E�s�?e�����S��T��'���Z:�v�:��{˹O[;L킡�
v__@f�)3@��P/�T*�_�H��������0����MC��J�QCg;�A��j;��"(W���-XY=N�6���Ce�kI挍�S`����K]���8ehxy�v��/[qI66���T����7�4$�#bԹ����ȋ0C����x�AQE�! �b�F���!�c�%���)��X	V�x���d-B�I0(��<��5�L�Vi�.��m����ءQD�0EH��Q$�a�wDb�������$*_��t"����^Af��#{�Fa�!��ɋ��k���L���G8�^��`s���E��M�v����B�r�}��2��\��y��~ԇw}Ћ�XB�	�����|��8� ��L1QC��դ��5��'[�HT;�/���q�[��{�
k�d$8=���x��!��d��ihڬ$��Hv����LQ�z��.�]�����RhHv
�8cZ1��8m'S.7$�;�>��-!�Θ0���.혿v����лH�Q��{!P�z���Mئ�P�*E���%����B��@�(�6d��@c�!�h&g�㎞0G%F��v��!��+hr��SP �����L��j��
�Y�E�w�f�,�fB@�Q��|�=��F?F�M��c���9��B��CqIF�|�r�
����P������'a���+�����~���jB�{���_���)�%Y��