BZh91AY&SY�PWx :_�Py��g������`{��t��;}�\ժ�f�C�A�ɓ&F�L�LI#��FC@F��2  EOS�z�4� hd  MQ5���#�z�
d�4h 2hQ�I��(�ɴ�m@d h� �! ��'�<&���� ��4�4�:���� ����>�q)@�>!���R�`"�V
0?�%&%QK�Dz!�ĩ)i%���a�u��mJ)N��"�,�H(Q p������f	�1�HAH������dq�3;���#,�����D55��d^L0��!�l���u尾�0�5R�	�Ǖ[���kYK�3l���K_� �k��%�N^�♥��ES.*7�f�3A�A�ٴ-�����)V�a u���+I��PB�)R������\�]��s�
��A��%���&��e/�� ���[C�p�v�L[�Q)�2B��6�aEs.!�	�#J壛W]d����J�c�G=&�gR��ʼ���{���F4��I(w��l�*".�� et�d���A�����l�lZ�9:<D;Αb(��U���M:M���FO�&zp�bЖ������Hh�Ճ��Y����Mp�$"��[�ZI�M�JRb& ��P톥�C0�%�,�����Օ�+R���S��x��&!S�R
�	`I(����@�D`j|����֗'�8~����)�`8Jo���g\�d�l<\|{�4n|u;��ϮN��K][T�b=p	��UC@:� ��J~BE��ҙ�M`d� �H5�'��A�̓���G8�W����LGv�|��O<��*u�`�!���9� �1X
�hI��ԁt��Lw )�IEFg2C�̧���a~1H2�)}�w��Ɍ:4	���T�$�P݇��c�r�7R�L�J��h(�v�Y���mqj2TywQn7g��ksXR�$���� 3��9�2�5��f�@��j3�|G?BdTKo��}L;� ��Dby8X`�����H�^G ��څ��e���Q�+<C�	��
���s��.��@X��v�񎱝H����LG�&�s@�F�K��3���;���c��t'�.�,�O�8�@�e��B�LW�'�;�f+���6J�X	]б&`Q��e	�����|�!��a���p��тY�F ���V@�K҈�@S	UA�B�KU���p��V�@��8=��ME�N�n3�I���'�&�A��2lڹ�F1�'������H&��j	���^������XT���)�>K�ǀ��p��vǠ{�:�NB���&师H*gc#�A,WS�uJu�q
��G^+:&��u!x*����/!#r�Z��[[�!y�T��4�X�݉ca�P1!$�K䠶r6�.��hm����RO!S�U�� ���+��f�V�Qע]�]��~��׍���A� �;���-�2��b���"�(HY(+� 