BZh91AY&SY��� �_�Py��g������`~���of�� 6=���f�P�<�ȞI�M   h  �4���i�@�2  �A�ɓ&F�L�LMDD�5�OS��4  �E$�~��� ڀ    D�j2dhF����zQ���4Ph��IvتPB� Q� �����2Ȩ��A������
�\�'p���B,�NQ�ї�������Ƶ�32�����3+331��4�,�`�~�v��ܷM���7S�����U���c��H]�Q��B± )_
�()���D�9���5������=o���Ƃ�'��2��]o�4���fm)�Z�t�Y��8�"W�6�B��T�W�C��z+N!!Uʍ!Hb6U��bT�Y���绫���X^s!J���hT-�������˳ ڐ�߫��=9�7*+�ߌ,�ijy��+�uuI�\rx�j�x�1uc��8�U ��f�ۉ��0EO��6F\+�u9"(�#P5a�Լ(�kZ!�G�� ��-��z�h��4)���RNPEC!ȱ�(�ƶ7ro�Y�K�M2�6���YۋQ�E|���<:�Pm�Z\�[������zЀ�/��Qj�!e[D ��������;��z�+�]GN�ܷD�Hkw��X�C퍇:�+�B�m��D�˛�$5��٨�f�*]�.��}l�D��h��e�k��ffe�x�II�5�l��D�ؤm��UѾ2�W#!���l,�
�7��r��m�j�`�^B�`N��b�x��Z��i���b��6�J�V��tM��ƙ!�4�8m�`��Q.�q�Y�f>�fNƃ4���6�?rf�:�) 2Tp7e�0�z�z_g���!�KsMk@8y�*�d0z��Hz�0��6$.�;9u�)�WQj֖��u�ߢ9������6�VH4')�	La��+4�]d2�A��+��9�ҚZ�i3tZ���0�
���x֛j��I%&�2\%��e���i�&"$�dA.�F�6%b�H��FMR~��Y˜]��M���J�E�Qf�8+����=~Μ���F�YA���Ч?���&����NOe��{N��~� ���L�<���zq��˧T��ד�Ȝ�:B���������#�
[L�2J�@|�${�#��&��T7�$�	ҏ�BB7�qY�a��Ʒ����[����]O}�~Dd$��4�K�^	���ۜAB�D���@����"Dy�K�ӊ�ki�+T�j9o��Z�ΌeZNюm�ȆE����D�%V���e$/��nkT��)��5%���L;fSY5UD�(j�6*�֘f��R+�v���{��a�H�7*%0r�B?����V��e�[E#�oO�L�`�⋇�X����J���y	�j��	�L�$�؛��dTmZ�2

J�ƋjY	`��L�� �e��_H쬫j�)NHl�K�Ih7�Pf`Q:|t�!3�M�!$��1��q��{�u��l ]����1�E��P ���KXs��WTSr�)�V	�A�@�#�!M 4f�0L�H�}e�a��!D�2i:x�Y$�nF�q�&���de����?O���37��"�(�y���>��{����y
��Y�	z�A�+u�G�qʤ"��ȯ�߇,���֊��ni:��R�$7)X�5cP�5&���@��PԨ�/��A���h�u�S�a��Y��\1[|n�L	��k,u��9�j���yx�%t
$E�Fː6�~,�f�0H����L��{CH�!����z� ���0H��8Gm)��zʶej1�٢6�G��&�0�"��.�p�!��Z