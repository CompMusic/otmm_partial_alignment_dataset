BZh91AY&SYh�� ߀Px��g������`�{suu�� m50���$�Ѩ��FM&ODш�i�h�&��@LQT2�@�   i��&�&	��0`��$҄J4��d0 0��昙2h�`��` ���DB�jm4M�?E6"�z��x���/D��"��HP�����R�H�@�2���ԕ>�I�@\�����Qs��X�mmUaÌь�6��JR��fffn����䪪���ŵ�1n�B��K7x��w�,�[�5z���F��!Ȧ�s���y��ڗ$	�m�7�0�,�Rh���/\�^\�>S�����tM9�];Զ����2��
�q����1�sI�
��*Lk֕W�u  �/7��3�M����u^��SY��iMa'F���:�(I��9QW9��U,�թK�R�&�c{���u�y�G��ɭC+X���J��r�3���&���BմDRJ9ni4����[+z$H��{9�R|�ϡS�J�f\�b�Q�wl��ۂl�lH�tϛp��s�,��V��Նp��Nj�J����3�T�3 TF ʱ$��R�n�;�1�k�^m���Q6���mEk%���ٲ	���a�ή��zW�����jd2aQ��7��W��8dԲr�jB
�@�v@�5OW�T�9*�$MD5o�&�E�K�	��%Oq�]�c��!�Y��W6qW_��D.
�#�]��|D��ؽ����	��#�4�U�Ã��f"aF�K��E�
�<��k����lT\N����T��E���x�%��ku.&)���JU���X*L�p+��f���e*c:������//�)��-�A��c��亙N��٪C;�����L�ˍ�iQi��'xhF�ö���Q� G]U�*�f��9�Ѳ"{�rzl!�N�V�jVH�R'{AV�K'Z9O-�p5� OR�Ƭ�3���Z�eZ��#ߔ���N�͸���vTE�*��&�.��CM{�V�U�����`�e`\5�flaZZVC|cxl���DQR���K�1�`T�U*Rؚ� (�ʛ��j�͜1d0���̹�57�P�3\��i�a���8�T�XaØ�v�'��ݼE�'&z���&���r��hz�'�ѭEv\w[�"���N����;=���ٳq�t��D@���?�B�x���-/�ڡ�%֐,��&ď" pVc{\�.�Χu���k��+��Q��=�f_��n�:��꨾jvz�2���Ei�TP��r���/My1��g+��oLς��8��[�� Y��6Z79�	�s��3G�T�"������7�EX��Xt������St"�tzu�tU/"�������׹cB8P ����C5��mj����rQ����W$��G-�&�'�3��r���F�+�v�0��`F�DG�>�E\76T��;��H�\�Qy53g�hu+Zf��T��H��z�/[A�j}��.�Z���S�ٞ�,d�'�u��b������ Z��!q�7+p�5���+ЍM��vԗ�A9ؒ\� ��Y������ y��/T�X)Ve�0�wY�'igȪ�F�9}�8�k�F���	�v�abHN`�����:�.�p�Žc�ԕ�������Ǘ��r����Z����* V���-�|�ۅ� �uYgE�D���@9�����畱N��W�V�N�8&����Nl�h)�1�Ȃ��2a��"�!ў岮��C& PVp�B�E��Y#G���14�{'��ph���A�@�ĚՔ� Y��	yvw
Y��lU��c�Ƽ\j�>��Y�"��rE8P�h��