BZh91AY&SY�+?( m_�Px���g������`�,���w^Ƞ �����n���R��Dɡ40F��F�4���i� ShH�� �     �I��C�4�44 �  4 $ԚMz�CL�4h  �d0ڑ�iOSb��hh  �� "H�����h�ڞ������#����pW*�7�%��3
 ����$���Ơ{�< ��*����p3 .pI�����^;wB�m�L�1)O&���y�5wqu+UT�Wwqv�x��A�QU���s&�Y�]t���vh`zg^3��3�1z)�з��.�Ԑ��ڮ1��L@@��T�j��-$�B@=�uA�uE&��]�;N&�!���j��)����eJ���ٓL�*#\`6K֔V2��|��y�`�k�z���x^=��<�$Ӏ��U*S��b0ɚ��-ramf۩R�Ӳ������<�LB�,��,���Wpi��&K�L�/�b�*��0�uX��]��P� D̎+�޶� �� ���:Q�;���8�E1����T8��s���pg4�/=&�M�Y�Rv��ux�4NS��;3E��'[��Ԓ�m6���ח�exƮ-B�rn��DAKCZ����fx��X��]��\���1݄RK�i	�!qeb�b��EqIn@uA�';2S���A��xɛ������G-���wk�*;H��;*�lm�&H���k|�\���(��	l1 U������D=	;ߐ��rOa]�c"S���/�̽���85��ۉ��.��Al��Ue�	�×�/<�/ևj��l Wׅ�t�ňy�Ӥ�A4e���*�d*��E�[-.2�st�����Sa�9���7(-�H6��;��o:Z�#P8��/��hCq�l�2:!Y7j;��wSw�N��L�s���B>ֆ������%)Ǵ�ĺ�kQ��Xd�X�$d����[f��(�4��6�&�Ά�ܾ&�#�����/1�r�+1����4@�E{UU	����C��J�?�2d�k#��b�JduL�-0�U&�RvyK��xaL�q��m!Au��B�EP�H�R����Ub�[F�P�vp.v���=dCl������N�W\5:[�e�.J�oYM�"��^^��z*y�����Ɂ�o�T�T]	�ǃ���4j��I�/]�����]��|m�b��sM�VD��;���sr�=L��>~�*<�O��Π2�V�YW$���8��gS�f��"4�U��	@b]e��
r,��H��m�Ǽ��5~�!>�������8޴E���������T�,�M*1E ��&Ɣ���H��e��O����C'xJl~#�Id'� ��N�S����'?yr#���oV
��P�f�m#1��@��G�Ȥ�_��^6>�n( na��=^�(��t4)��^BuK�q�L,�5)�w�DK�$�5�d3f��"�Q�8P����.`���'f��}�矮=z�]&؊�7�=�o�O/QيUD����8�EG���y�)��� ].V�0�@��&E�Y�
�X�,&x:�ıbQUQd'�SC�7����ў���q��v���-<T$6h�A8�K�P� "�����ι��Y��L�sf�k���[�p.��>�9�͠?��=3�t�<ʍ���aўGnY��rN��FIu�_YA)=�5ݗ�c����P��Ǝ�v|!`YT�%��#b���m3ْ���MUIVо�G$�C�pב��N���Fݕ�����X)����������I�ymIgdKYH	X�h67�A�}�'���2�B?�o!�V���oZ)��]��BBЬ��