BZh91AY&SY���� E߀Py���������`���7��  �'�����;;�IS
h�#Oj&��d��hM��S�JhP  �#    s F	�0M`�L$�E5L��hѓ'�Pi���4 ���"OSi42z�?T P �C �H
=#4��zM�h���h  �� ��o"PLB�~�bTZ(7���=.�U�������o .�UuEV��;�4�Jr�5k�Vr������̶��������Y�l���������x��hIפ=/E@�o��F���xS;U��o`ѵ݉�i�civd�(PB��EYQոܥѬִ�f:�=/2� �q�u�z&�?Q����hD&^����JG�\�n�)��3Ksծ5֦t@y\<�"b���N����bA�U�e��R�k�9�މx���Oc�����r�7Y"����K��=:�`�00Ds�|o�h��j5�μ;�I=���Ą�y	��鋶-틼X	��"7�ʶQ�6,�>^�CWT��"8D�mq�ZP¼��;J����9�㮻�p��`�@��C-�4�KU9��\�] q]�8���&��)9=B��Zs��c��-�P�/k��/z���Y㎶S��,�����6g#.�J���:�qi���f��b96�e�Q���3ip�8C�hS ���p��tF��p�CCtR�i}�qѕ%�������!����
.tA��k�����jl\m��P�����Ԉ�)��	�;�	�*v��yT(t�MJc����q}�	�UD�"g�X#�7��~��o��cȽ@����	@�c�}D��I�&�쟡|bG6c��秗������&QL�'b����|�ou��d&�ktk�E�r�՛����(8�K1҇P�=4Sb��P�Gq��g�n�<��y:"�!2�v��Q��0[��kD@%x���Mz�EWv�D>i�S��_9q����89������-��B�L#z�>��֐ ��b[���)��g7��g.�#��(��a�=���|}�c;mz��Bnc�S��V�\�ܶ�-�4UmQB�l�̥HT�[h
,�cpU�7�+-mU��E�CTX7�%t&"��e��[QK���P�%sK-��mcdp�`F��ƃ"��0V��C����R��,i�P(�\:%O��a�cS�ܞ��*/�=�MF�l�0�� ���~V�v5�g�p��t��X$.�O:�S*�-L#��%���1�DBE~�FE��=4e*�ݰ6���(৷ G���4�h�����=}�Zp0�O��&��Я���;^�]�(���S���u��;���p��j�l�E�z\���g���J���,DR,X*#6!'}�H{���P���eI�%Ce��'|�1��#�LBHDJDi	xL�o>��V8��R�S`�'|�Z@��n%aPK���7|z\�SH|�.��hEF��OEa��"u`W�vǺ�
?��c ��)������-�8�+U-�:�J�Ұ����
�d�ת�ݼ����2��b�3J�g���&��$���;���jz��v��ixԐ,w`�>g�-�@����T@e�#e�n��0�,�Eza 읾,��ν��	���0y�����;e�4��4n���l���Bo]����0�Ò�vh�3�<f�%��z2�PZ@?�{�[�7R`�PIs�Yn��a�G	kdF�SQ��"3�W ЈnwyS��,k:���K�r_��`5.@پ9�� VzW��bf4Z>.���P�$;g�������ֆjaY!��E=��;wɂ�PX��3�%���Y�A�8�*��<8X������'�
�:4Ν�outGQބ�G��۝��MchW��Qqo���tF��:�� }N.�������C��U)���U|���"�(HO�ZK�