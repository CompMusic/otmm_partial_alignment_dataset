BZh91AY&SYl0� �߀Px��g������`��w�zs� �>=�wvV��a$���FS L���4?T<�@z�hz �@	@ �   ���2      M(��@ 2�    I4���)�g�&�4� $He3E< d �M 4����Uk��`&��B�b IX��I�d؛m�jv���0@����8(e��cg�D�a	�k�ηm���J32��ffffde�5�����̍�C(X���i�w-��5�K��Ae��pU�!��B�VK1[T�iҖ�p D)4!���?n�wp����R�,�̝��NCO12���hŢF�!����H�5���Jb��K&Y��n&4�3���F��\�'"�%���Q�H
)� UgEQpMh̶�I����r�gs�Z�4hύBνv��/.�q�"9I6�	@c�*Ȓ��NQ����YI�!"�0�F�Ue	���4#����w�0�q;T둩����U��lr�R�@x�
=$<�.:g���th�B|D�@3*)!(������z)D#���i2l�$�.@�T�1�a���T��Q�q��JL�6�ɶ��u��qh`˪V�����SIR�b���E���^bC�c�zǘ�A ���-���S��#x��XVfC��^:���~wd f��m8��@�P?S��*7X4�����l�S�Ȩfxv@iW
F��i#�8��J0J(imH�FBs�����5��F�����jj�h�jw8�Q�����LX�4֡�������a�SY��rV0�	~e�q4�F8E��a*���F�F��ƛ���}�l���9.ʣR�����n�fCR��V�m}$��6j�C��2�
.{�s���^���#&�f�@���|��|t�`��g��:A\iVt[Co}�qd.�9�1�F�(Kc�kz[�YB�˳+t���e!�pޭ)�2�V҇Zi��x�nv5ǀ�QW���2R��_��8<�_�4�HH����wYQEFp�X�rB�V�����b��)�A�3u�a�X�`7A�3.,V�I�V�d�X��Q��S"l�UE���ܱQE�R��;,�fo���a��fug�a0�f(e':�����>��짅�`�>��y�'<a=�5��͖8�,�ϫ�))����w�u�WFZ�[s�wSpOz����棟7��\���K��C�.		p#�� Cb� p,OHس��u'"!$$��B/�;�A�c��t<�-��SoeW�A�ZQ�$[Tc�7��5����zgm�{�箹�	�<�IF"���^�w�h�ņ�T��Û��VI5EYm�ci����F��2P�烊�̜�|�% �_�2��0T�]�HQ/)`��S4+e"��p1�zF�aؐY9���B_���1>�ݍ BR��i��A^�h�R���P��Ө�̳CY�@X�#&wz3i"eZ&5��\,ukY,��%�BU��HI�ħ����Տ�}4ӥ��[��3��@����_h�*I�)l(���U�h�#9���dgd^6H��P�2�b@g5����zI���!�1� E�D��lii��
���)[�K,��f#!A	2d97t\	��F�	n�&���$���u�Sv��X���nsV[��6u����!���m2Ql� `�^�	�"��Jg�����<yCP�EVTU��0��@J�p>�.�9.Uf�v;�/��(�8BXXۦ�ά�H��-���dD+�XVD�+����{l��6�����|��V��Αo�Y��_f8
�4��!�\�B��J�]Z�!)�@rO��o5�Y�Tc_X�3�:d%p(��Q���)�a� �