BZh91AY&SYM� ߀Px��g������`_1�e  �*�1j�܄��Sh�'�{H�M6������S 4�jh4�H��2h   �����F@�ɐ L��  3ID�ҚG��L�bd`&�F	�i��&�&	��0`��"P��h
���ziM��� �hz��1l����,�%�2�Eg��Q��h2H�`�i�Y�?ͅ)<� "$��)��<g���x}_�����8��ww�����uf�l�VV>��!��oػڏp�����Ӈ*�2Xa�0O&KL�uR��_fL�i欪����k��ؤ�9Yxb�}&3��I>��!~Y��Ý�q�5�Rerd�QE���E�V3��Δ37�F@"VU8	*͛]�%Ko����ƺ���)}�BRctR�y�R-��!Z4�����x�������/�	'"Wzm���7��.SZȫ"R��c�Q|`(v,H(UKK��!&��涙贾�!�RL];8��辊L���-*Q7!�Q*a�/-���LL*0�A���87CKma��v�\Kj7-L�J�HBi
PA
�DY��%V+�L�$l��ccPĵ�y����f�,��
$<��xq-�<U��QR���$�`�H$�ń$�a��URЄ�r���̐%R!���xE�b�n��,�q8�P	�V0Խ�NF��T�D.�N>���wz�y�	$�7WQA]�G]��3���SS�4Pn���Beť �Cd��Z[x�bN�Zdd���}��ǶKXUy�ɶס�=)�O�&bqh�G��οl�
��5%RYޮHV�P�"��VO*���Ec��ͯK,���6?&' t��uZT��l��J�~f���
� 
��uz���f� �����N�=���}�uٗ��wi��+�."^rc\���氭D���V�6X��T��P��Ł���P��b��:X����] �@Li�[��}jO���+U]Z�&�*�E� ZFbFB� ab��BQ )�.(�F��ig�Z�6�����S@�,5�&`�$����ad��W<�9��AY�@�V�n���m�-�J�?U�ڠn\m���!�U�w��6\���x�Z�Ⱥm�ϐq|�[��rb��I�P��]�]kj������8j]B���EȠ���5����U��ʒ&�`�������%ĺA
�����f����T�Jb�=<G��a��KVr����T3[�� Hm ԥ��`\i�J�sP�JM��z��4�q���aIA!�)BA����CS�Ki��/Z���T�g|�F�%���F��v�h���caK�{�Y8�q!����$�`���s�*��k�ZN?R�)��'��xVj"�;�̎J���b�6א�o��� �K��8II�-/�<Ie,)�cs�Z��G���!X��Ba�Q���6��ϟ>o����
�7�E��~bq�g.��0s� ���ɬ��M�TDq�M���%uL�9�t�W~ZT0{m��sd
E-�"� �O��e�By�x�,�n7n�84�hp��`9v�\I�jn{x�A����s�oW������˕���5���O�6s��Olm�s;"9� ��Ѓ�Ϣb\��@�㰖�+����mT"*>Ez$��]J%P��OL|ĺ9���F��He>g��aE��E��T+�'�,��3��z��3,��6./���(v[f���_�5u@������v����2u;tQ�l��ᶇu�'��axe�B?��Vct="�}�~O���)�h^�h