BZh91AY&SY�� �߀Px��g������`�{q��۴H:TJ@�� j��6M'���i1����EM�   @ �12dф�14�&���I4�F����Fѓi�h= sLL�4a0LM0	�C`FD'���?Jz�MA� dM=F����u��TK�)�(jP
 �_�O�1)T
�*��v��� ����`f��\�:�v;�q��k7_;��Z�33333332��ffd�ٻ��}ne�(_Գ��j*��z0��y�ԉ馡��=��%V�-�N��$����֤��������#�2��9����B-�q�� �@�LX�k�;|	A�����U�.���I2�Bcf�$d\YXסn�<�`�)��j����tӏ#����rU-;kg�g���$�MM��ȓN��,Z��3l)g�G��O�p��C��*�a��suz:���Ưc|.8VՍ�u0�T��д�	\��4����=��`��q��p��t�"˲�\���%z~.�uB���|�#�tnp!�H�ɬA������aAЕ��Q�@��qҠr���G �)��5�� aH���Lp3]�nq�ӵ̴Y��b��]�l����h�w��rj���d�!x�� �\"qfIK��֚��q�f:����+�[9m%jJ>�q%$�9����l�u}�� ��s�:)���@Y��J�6X�Wf.@QJ�(FB{�h�����٢F�#0�3J���jS��C��u�����ZZd��{#�TX��C����]VVъ��ާ`�Ye�Q��Ԝ!pc\���c����;���ӈ�f�["�ĝ�n�> =�F!O�C�*�dU�)�R],`h<�vMW����圑s�	�!/�8�t5�mg��W�
VD+	H�Ӽultb��p;�HX/�c���Ej�GH����.˶˱q�IP	eB��O� v�)�.N�@�n����+�6�m�֝ո�\�d������W��mup�(K.X3�9�T�:U��WLH��w�VV)"����v����QW�UPh*�'[>����G�⩨��A�
�K���p�0�A`��3,��C��-Z�EE��U�� ��G��(Ҵ*�o��*�##KB�ѵ�
)�!HՎ�F������*����M�)�k�.e�c��̐&b�U|"m���ڝ����V�{ԏ�~3���a�N��,�)6�f^;~�:�Y��Q�#��}6��R�u�9����@����}/WOxl?|_��Ծ.���H*E ����m�#nܦ�Й����K� ��zl<��9.���UѤ�^���b�=�s� ���xITR�q$�!�o�wx�h����6�e��Y@���ij?&��D#�/$˅���6^��U)Aj��Z�)JNb��S!c�C���YC(^�~�&A�?�A��E��i�o��q�ѣ�~��������䆕2,%`	l�_v�E����iI�❚&�pd	A���%���Μ�uoR�TM���)Z��{���R��o��p(^`e�8f|����Um,@������o~$t�}��e�hl�͌�IL�_�%�#v�a�P�Q��;�X�|�:6)�R�Dt��2a��ɯ�9� &l��	��i,%�X����(��H��ӯ"����e���>85���+Q�
����ݘ3��s �z���v�h�����0��T�9.h:�����~���� ��:��s8�@��`�N0�Ϣ7��@��%3��Sv�޼��v�@n��錌��<JT�%q��O%6��3�F�*��j�0V(,i(kn��kW[���UZ)
3�K�x�_L�7��Fʋ[6�ެ����99��͟1c�4�\C��10�xm3Ax].����A�sl��:\2�x���W)��;��܃l��w$S�	
1?! 