BZh91AY&SYEv� �߀Px��g������`α��=�� ���	��BH��	0�f�#�hڙ<SM�i�A��)C@      �<�S��� �     i"�Q�����d�  =@sLL�4a0LM0	�C`F"@�&���2z��M���22 l�тIN�9RB �&BAB@ �<G]����@�"V�>`?� �@^摦`f]�vZ�4�-y�l���<5k�cb���n��.����ff^fe���B�~�ܧ�7B�+�k�D0�&eQ��aZ����:Z���Uڦ6�H�%�+P�w��p�e�7��Ϯ��u7���	hh�������P��BU"���4޳YQ"�(ڮ�f*-�,�WhX[ը�P"4�,Rضa�)���V,O��8�p�V�ŷ��5,U���`%I��*��	4����K��%�h�Z�7� 4`3 �h"j�#��L�Lq1T��}��Pӳ6���� "@&�ψ5�$�a�M#Bw!ck�ڂ�ȥ��X��PQSS����@Q
&u-�X�qW/q8C3��NFaΰ嚏y�z�s�p3�3��D��(@q���b2i-Q8�|�!ceߍ�|,*:��+�`�,E�<5(6@�ei�o�(ˬ��|���23u" c�D4��*���)dQ��x�H ��:]�ckX3 Y_xm��4��I"IRg����m1���H!�F�����9%6��Ŭ�5"K�E4��.���QK˴
P(��Ñ YI`��Z,��Ȏ:x#��f�t�\M�`��h۴+�L�8��m�i(,����W �"��|a���-f\f���	H���ćM|�����a�����WzTB���O9����+B����VR!� h��N	��&	e��	� t\��	Ѭ���/r&�y�ʝ�.�4 ���z�'��u�[/Oׄ���J�wj8y�
8�Y�ඤ�W���Ǣ�ɾ>	���$)�.e%�q!�(����:��=y{/'L�kw���Ǝ�vO)쨊+骪	'gg�y<�1����ٰ��v����UMӵ��a�u�l��L��)��&�b�T[^-�1�U�����]2��e�eeF���8ɉ�U"�Q�ؘ����-��q%@��q�<�6��bk���bM�!����G��=��������S;�0�G��1��hz'1���[�;ry�G��53<`yu��,R�=I�� �-ܟm�=���\7��X���!�/ p�#��o/�e֞�B6�$���^c�u��ط�+��5\+b����ʢ&�:�(!l^���&�PC�`��G�~�'���[`�P�ݮ����F�>���s|(iHxX
��Q`�Q�Yl���@c�[�p��ׂP����6S,�Cc!��_Y���&�[��r@|/�41 ,j������2��iW�_f��&P�p��[�Z%��̠7FBY�_��J,2Бu��#D�9Q!AI]�}OV���ف\S�6@���y��I'6:(�����)[$�Ys ����#&s�d@��E�9��K�r[K#$��� K*�lddږSK6^�5/>ɐ��{�����'�CD;�q2tOb%�9��I�L�v(Nl���'�}�����!$��ۧ�N �
ԃa���n�7Hb`[G>V��5����%�H��
��J<�%�(S=���W�G�u����m4cF��ԍ ���^�`�]m+���)�1rF9�)P� %LwDF�$�Wpt�	^�czfk�vPVXA �Ye�F�7�LM_�~�GXKU�A��OU��%��4	H���<�G�ܩfaQ�1�gdO�h!�Q%���.�p� .���