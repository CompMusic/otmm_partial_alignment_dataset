BZh91AY&SY9� ߀Px���������`�}���s� y�n���	$# �SMS�Љ�1=@�4�I(hdd�  4  ѓ �`A��2`�S҂Ja�SCCF�    ���S#M&=4i�P�ɧ�M	�4�����)6Sh` k޸��O�ڂV�%�!���e�s¸2H���������w2V�lI*�r�q}y�{xq���|9^���zf[]���f>ffFfcb����$;����b� ��:΁szpxJ�4��]Q��+�qw6���N�u� CYi��R rR���c�r�߉o��͌�o���71��Msam�B�[�5�
]/iq�)Rdަ�`�iMmG�������3\kĹ�UՙS���5װ�������q(/�*	F�R�A�䵖��с��0�4��r┲M���_�^V-6ۙh:�dU�7TQ�J�z��%��n����d�eq����	���ഃ��[��.��:�zC0��FFr/�Ѫ;-�OS��O��hB/j�L㘠	vb�#6�� ���4�&Q��ʻ�>ဪ�^� <B�ј��q&�\��� ���W܃,�DR�k.!QH����.�OJ nѷ#M ��o-��!,�(���m<�tVbvB����D�R��ܛ}`���_	�͛��EY��fh�((�@��:&��˄Y��'@r_B�#=��ӗ�]X~^������rD��tn���(���@��#�V ����~jƊ�޺(����
\M68b�eVk4��\�r���\�F4~Rm`m+R8[Dat�M���pA��8�]��T�(�dҺ;��*)� ��J�@@��
�z�^z]�_B��ޏ]"B�AJ����΃ę��� �|i��4N�e��j�Xy���"8)�0�'8�H`��V�+"@,��t�E֪�4QL�����i����#�l��`q:��u���Hڡ{j�GT%�B#I�RB��U@Y%P��׌�#�k@���2%�U ���bF�	H�N[�U�D��P!��XѮ<]y4Paf�,�B M�5x�T�������S��[�u('�Qo�O�#�������S5���ƪ�m�]D�g��u5��z��Or�P��\:p�xFߝ�X��]kƈ�L8��H�B�J�g��`�a�R頙��<p��k_��1��� �����~�(b��&a�w��E!�Q��/ڷ���}n@�T�]�/�MJ��k���H����A#���:�*0���]���9��k*�@#B������Mh4�͔hR<H*9�⬳'8�(EC=���-`���������k%��8[+L��&�/���<"� �h��G#4zC�\����K~zSB��<9H,r6QХ~��z�Qc�Ӵ����G��60XƃqC#3n��j\K�N�]`��7�!1�V����~���_K,u����^�!'x��b��Nҥ����1/�櫰h�#q	khB�dmdbڑ�O�H�� l4�
Q�)�HE�$�D0Ѓ�
b't�SRf)�d�TE���+6h��	�£^�Il3��Bۤ���&�'0wuH;���ֵ�CdC����?�6�]č�S�q<*�~ y��˚:�
�@B���)�8ﺃx�J��V�ni3����9&�~[]zޱQ`��.J�|(�;��6QD�)�ӚV��a�AJ���MM����H2��^&��8�d�

J�H(�e�5vY#_��щ��(�8e�ʦA��ĉM��HB��\�'�n��m��<
�f����#��T��=��]��B@L �\