BZh91AY&SY�]ʱ Y߀Px���g������`�,Z�q� Ͻ��tn]�V�	"�M1OSL���j��S@z�� �@�$`      F%OT�i� �     	5$Ш�����6���   =@"��T�C�l�4hz��@ h"H������I�4� @dmO�4i��.u�ވ�@S%� (w~e?8^�
F5�i���W2 �,B�` ��V˳Q��/�Ì����+���J>e������e�Y��������՘�/�Y��	`�|a��]��)J�g���v�YW��Qad6��
b����l�Q>m_��f1�y_8&����m���c[�CQY���V���T��uط~�����+Bȉ"�ؼΞJ&��<���C1�030'�R(k�

�6��<܈�H]�X$E�Ѧ"ɓ۾Y�pN�&��u���ǢA6�գ��F��I�.fI�@PSR�a�Je���L�0d�RAr��(r�"�!-*>I�dy\*V�m��d�V�n�/�.�׫"9�bl�U�e�C3�1��;�!�U�����P
Im[�Ŵ�� �-�Q4"8��W�Q�C\p�05��:��n�3p�),~_9��%hp����m�Ռ2��8�qt+�K"S=\8$/H�� �
U �쑣^#��z4R�$<"��w�R�i��Jۈ��Q���H#�B�|3�uD�>�by���Y���ƋJK]qn\,�Y{[�C(��ND$t8w��V�E�qTE>Y��D���-M?���*�8ppi���]<AƇ�(h:�>#k�I�Se��``���<&wb�dֱt8"�4m�wfj\P�CX����C�%�)`&�d�~K��k3I���X�j�͓��`[��{0-�n�;
�U
;Ⳕ Ҧ�Ts�����$T��?�I�z_Ɵ�x�/����gm�1�p2����N4R`��mĲmm��c�0;.��+�fTz�teF�`���y�3�[&��;
"��*���	��m�p�m�zָ]$#W���ih� 6�I��E�N��b��
Qi1iYf�	d�b���-ʠ���`����P��bEͪ��Lmk�0B�d��f������0��L�t��`Bf+eG{�������+��v��D��/����ʏ�j���N��J:������V�l�Q<�_�Z�N�3+�N&J��V���6��6p_��1�F�r�E;�Pd�;����:>��k1d
1�m���c3Ϩ��s^��B�0>���M>r�+$��!�
x��K6�Mؾ~��hyU��B���vIU1!\v�2i���!gԛ{��eP�P"�Ł��܀]	|(pլS(^��VL��ÿ�8�Ld[�8�4�f(�x&\�3T�
�Rf�c[�^�$���$�,�6���v�z܍��	�
�t;H-Ў�~�ImQ���J�c'���4lH�k��y3�n"Yy!�f� �{ܷ��^�-�B�3d��l�L���C�T�9���Oa�$$��(�z_ 9��VIU����1�(��G �I�I�d���*%h����(�� jtR�	�-��r�1�T���)���re��F^�:�L��C�`O�W ���(��'C���k�*^w�P=����2�oA����^6��� ����H���MTt��80��pM ��s��0ۦgfz<�j�/"a#$�ç��gPg?WE��n�-�&�r����!��KK�1�<\��v�M��8n��*���h6�k2�)�(�BrPʸ	�l7I"��]�	�C���Ѝ�!�`���Z��6�5Q�)���ߝU�H�#k�P��V�
��<���v��ܑN$?Wr�@