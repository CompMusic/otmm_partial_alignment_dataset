BZh91AY&SY��%� _�Px���g������`~��3z�   nz��v���	$�0F��S�2f������L�D���C#F��4d���`F�b0L�`����M���4@  @"��S�5�� ɠ   4 $DCS$���~���`�j � z[e(,�٤��(���UY F>�O2a)T(�QMD>�����
�� .�M��%t@`�.c��_N��/ύ��Zֵ�]�|����������}Y��8�� ��e܏d�[����Ш���?�vj�ʗw�̬|�s��Ђ�1�.��ADP�b8��3�_�&��#󹝙��I�ݽ��4��5��A�6��!v�0)̎e�y5&ܕ;�z�Q|Ϊ	#Zڼ��X�ܥ�~S���0W+U���[2&Z
"Q9a2�B�UvN�ñyy� Bi�7�����nV���U���fA���ū6g1W��C�H1A�CH���A/����V�-Q3��Q���6�q֌i:��'bɟ=���)k3��������m�.��b	�,�.��� P3>�ۧu	3�1�DX@u�C�L�T���C�sL��L]̈�H!��/�$�
9+@��/�eN�D�63�@�Ȏ����5�� ���#��XA��O���e���n�vyqE���<��QF5
-����6A9p���Ɠ�Xr�i���pa��ݰ�@�m� i��rXx�����F����\����{-:��4W�]��$L�g���҇���Ed�=��$rr5ox���_���w�΂Z�8��Ex�:|6����ߓ�Psg���G-=� ��F�n�Y��|YP�+����fƨM�B���O��g��#�}�N(�ޱX����ǩ�GHDE�<f�e��,G�>���T���dk��T�'D�:��{�����ۂ�L����n����O�N ���^#��(��UA��`��:��D���S(�^A�Ṙ)�p�9 +jʅޗ9�5Be�jH��$*!T�U�/�Dr�p.]�&r���b"����eM"�p�$i͉���(��*�u��F�ֈ��1h�aF��46 �0j�V5�c{K��U�辿J�O;������Bw4:ӓ�4ab��w��:��N�.����b8j���ڟHB��/70AD�Y���Xt�$Fi��B�䀉*�fA�
�
��	������!gҿc;�4��.�m�n�*����62=�Q\�,�J.B񾤢����Bk��loz�x�D������a��8��	�{��o�aF��i��DAij�AQ����ЫC�N�������r�\��w�!hT�A��	\�_J�so0ⵝ%w�@��C(�Z��<'��B0B�P9ˬ;�ģD�8v�2�
d̐�(�|�¾+ϡ<m�\�f�~Xl8���'�����3�S�V�D�~p߄d�ξ�- �hBc�,���'=���Zݎ��!%�HJN@��޼ i��UZJP��
Y���#���x��KI+���i��jr�� �`��d0�zo�Q��h6X�H�-�W���W�)e�/���'t���T�F�4k�&�j..\ ��`�$���b�p�թ��9��l�<�o�N�<�2��HġV���Lb��F��P�B���+��/�v] j��H�i�D���@8R�~�M=�^�)�`g�ϣ����uQKw�J�4��6+&U0�DD�S��Hz1pk0	Z�j�1�Ř!AYۄ���z����yf�Ѕ�i'�'�P�7d*���Q���W=���F��Z̏������~�4�������,�b�H�
���