BZh91AY&SYݿc\ w_�Px��g������`�,Z�qB�7���`�J��$�=�z��d�L��� �R�L�4 �14�# P�	��4��F��F M4�f���F��P  ��&MLL`��D��$�
~$�)�S�i�@ ���k�+�z�
%��5 Ow�S�B�d�P<U�e����WB �1	��'p��Z�t��1ٷvQESKS�wwWv����Mb�������s@���c��]���	�J<u��i=`Z�$��!�Z�*X�
��y:	�K%�^" B���F@�x�\����wW($�������;�k�Brc�/DP�!kk�Fu�����Q2��HE�л�M�b��+i���2�e'x����^�\���,�b�3�&�Lÿkڨ�b3�����&�m�_��n�ҭ���XrT�
U�@�r�R�a8�-)++��j�UԔ�R�����(��$��ʥSA��n;4��ݚ� ;G��� ^e�o�f�^���+��e����a`6����p�����Nƶdkf2������������	A���s.�F����<��c�:@�M%"d�!y�RҼT�K`�!]�2�YN��[ʿ*A�nP�I\��0���R�������I�X�F����I�s0�LE�7��Z�
QNLq�	L^0ٛ�q�3C�k$�X��DاƁpk�"����yH��m@
/#<�/���.(�Dt��r�$��K��Ȱ�LE7&m�u0,Сˌm��#(�Y�Q��y���ćK�Z�ZJ<�&f`�cbZ��С��`�a��A�w��p��bӷ����D�&AgU�E�*��LXg���b��⣎ט�7�myp�|<��_UN��.���e`%����j�����������7�6pa*��2+!�m�������@���חO:�li����� @p  ��l�]�>ou҃��s�V�F�d�N*��A�f	�K�$jH���&����'�L"Z�O&rⱧ�(4��T�	�B��Q`J	U]ZD�q(3��8�<�p��Mq�|����������*;��H�Bn*�<�~Q���D��^��T��f;��ZY%F��(,���S����`�/���yC� � �ppRE=�(4w����n��2%�W�B�ּ�3�� 2jW�b��I
��p��#�VIG�!���ݶ�Kh�S�7��I�̿����P#2r��r�t{�`�L�����/f<�d�@ȄV;��$h@�$ 	��Й2�%g�{֘�f��]	��`�
��j[�t�]{���t���K�������S2��.�$/	�D��X��XD���L80	B����gm��=
��Dnh�U�n;I�t�$h���5�3�DŤ�E�,A�ױl)����B�30	0ؔ��e�XC~Z����]zA��̬��sJH]Z�0�����qfr*�`$��0R16)��� ]w+yV�B�͓��,^�@73����~��]ՐX�˒���Ȣ~t�Mk�,�l3�9�3}Xk+Ì�FTGgo~��I֨��.���q��>��� v3��X �bwj�y���p\�;�+@.���t��NJ�xaQLu�#�U��I�
�|���2fi�c^���L�6~m�z�AlT���N�6�#��[�\�8�����M^M�UU��x�f�mr��a`�n�W+�Օ�HNF� �]�f��.�kt2����Pm�K�!Ԩ��&f]oA�������~��88�dB>��C�z,� )B�Q���)����