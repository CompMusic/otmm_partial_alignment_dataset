BZh91AY&SYl�&� �߀Py���g������`�����o�����)+��nL�JE4��=�M&��y&�L�OD�A(� �h 0�� �A&��)�       I��I� `hM�3)� 	��R�MM��4z�jf�  4  $�5'�Si�4  	"�]��J�P
�܀VJ�>�nW"��>T�O�$�M�!�K�� V!]��F�0��q�g'.lc��;�����UU�yTI9Yf�0]�jN���܏l8s��.\���B�]���pA�$fS�7�����.b��H�n��IiWe�6��Z2"q���9���ޝ����,K#&O��pa�$;o����1�2��Z�#(gmц�`ޔk��2t^g~ف!��a(#2���#�^�0������.�6x���ީI����ju[�I�� Jr��P�#J�0�6o;:u/dN�b���Slu��cp��k�f��yX(�ׅb�X�&}v����e�4	�2�e��MY9�%��.o���׷�p��e��<_	HFa�`��!A2��� �tb焀Պ��cu����Hgw��Z�@$<e��D8��ө�.��i|�&��*�ޚ2݇slʳ���%aP
ۍU`��)�\<�!~ lD���J19Ҧ\�-g"Bb@�ա��:N��\��7��J=��)\���8���ErA3�L8�$��ai,1Bn*��bE��bXS�P!S��\�|�;g9��X3=J�(�	ZI�[����0�1�B��@�B̪�L7�5�)K_�6n�{��zO&)�Ъ��!4)d`�&C�ȫ˾�Dr���*�	�y�����f S��p�`4r/xKb�p��µ̲��Y*�1���.$q��TS�06��KEWSx�yܤ�i&w<��KO��,����tt�Ih���VF�k�!�U*m�&��uvn,/LG�O�:�H@��e)�[ �oA!pts�"�ٶRZ�&&n�cr��1��Gq��v�	3v�%�X�'��KRdj�%\�[����mFq��\�CiX��Y��N�r*"���PHHП��qJגey�����sT�mB��e�M4%<�A�
HRP0�Kdif�,��7b�T�&rk�A`�RȰ-*��-�"%�Ћ0�ej͔�Q�4Pa��7!&��vaވޝ���uINlt�����x~�?Юhu'PzKN���I8��������>)'��\��nQ@�Z��t,u��k.����6[iz�sL�7�QDA���ʝ���
�̱�/�-�j�ؗ5���]��/5y:yA��"S.� �RppX��{җW�"�"���%����W�R�)��"�8Yj,QT\)P�*�N�@�;P��e�h�r��,�4	t �M�Э��鬕��gV6	�rzF��H-�t	��%�0��xCUq��W����ҍ�ܓ��l8�Zˡ��J�m(/m��#/(�����Uz�[�h�d�0+�%HN�a�7���PE�^��|���g�=N����[�.q2.�z�N�AL���^'�j�
X:9� �#6�dhb �;,���+nV	�4URBOM����ù5N<��M�dP�E$�,��%�,����-u�My$�E%/��ޕ���ViK�fj�u�=#��Q�,�-:�� ��4���$��t�p�&9�q�KʹgE�ni3^��&q��ͭ���2_?�*��"�ʈiR'L�a�U;�z��K�@j��ȰH6es�8�a�J
F�ȘU-�jߪ��BZD%�N��f��2vKm��A�15�F	WA	Df��8d�~�Y��ƾQ�3�;�H�"5���w$S�	�ip