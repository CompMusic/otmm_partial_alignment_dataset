BZh91AY&SY3x� �_�Px��g������`���N{�zM     =�!��P�Bhi��MQ��h	�di�4�mM=Jh"������40�4�OL��=A�@     I��P � L # !��`LsLL�4a0LM0	�C`F" �i�L*z��	4�z� ���P �� C�"
� �i�ϳ�� d O��'���`��Sr؄���\�8��������?���L:i��i��i��i���izi�sE�4�G�i��Ŧ��i���M8i�w~��h�����+�>/���ýT���Quֲ.��8�sh�Ci��TL���qwJr޷�[�/ˇ�3SSZ�#�.�UR�QR�]��)#��	T\q�q��[�۷j�tŶ�����5U��I�MT**�}���K�4���S �u��Z�&ѭ�*�4��Z�%��e���r(��R)(m�)3	QW�����*��)A0�2�*�����l��/�bڮ{��WL�A�I6�;(MI�K�շk�=�1�X����ll��n;��� ��9�͒�*QY��_�GD c~���9@7*�F�"Ʋ婝����)�#j(N�0�(G��UwB�P뼙��N��L�B�R�.�<�V �b(�i'���E���q"��4f
a��7�l�a�$�'f\��ac f7N�DbgJ��K���P�[h֛�/F�s�w>���D��e�M���!��?�~@NS$Bn뵘�۳�T�3�	6�ś�vs�K �ǋ�z�{T8�ut�s5�z�]��س��;��5�1����gM�q�$h��d,�S�����u�v�Lv�u8�;�S�j�ä�#�D6bC�xCN�qR�v�^<Q�K"�[����J�I�bf��������$P�,�r���D]Vk�e{�_���-�1{���b��G"��/q�a�\g�mfG��ƛ>��WV�+6;	�G��4�r+�,���2�=�E�g	����zN�N&F�q)y)��Z��MS����Q�����H�Ad��ۤ�����/W�f-�����$�O ��>E�D$�]kUWQ��Ҋ���e���]�&h�?��zk�='����Fy��J3��ҘtX�|=�׺��zG�"WQz��nv�.���k*�l�a�Y���O����8Y�s|K��Q�X����Q/���Fd��iM�Z c�!�%��]V0��I�裑�,�{t��y1i��_���Su��g�<c�!}��T>�3��!�Lh����:��EqpDl�!#�'�'.!m�;ٰy���we.p��/�x��;F�\��T�Yj����]���ȳcf�4֣1���iwc� �A�+�(Xq��	�v�>\v�&�O	���܃w�,�Ȟ-� �������a_�Oɞߔv��WI��ӣ�C�����1ʢ5F���m4񇏆�N�� ��` ��Bzqɇyvw���Ou��o	�}n�q3�wl�e�ͫ����!��M�~3����:t�A1$?v�|r̓�N����tόX���lKq��qC�Q�u���8]�H�?��A6��Yӄ�|`৞Ý}$ޜ�Α u�)ƃ	2��_:������Kݰ�6dL�ے������ӛ��j�đ�l���֯+�Ë�ѳ����8x���E�*�d י��y��Ef>u��V��M��݌S��E*
d�D�54�
�D�E$DvpLb)'}�ޖ�����.�`J0DL��dAb���M�	��d��DK����)B4�����#0%Z5�Ѵ�)KJP���C�"�	R%)D�30h��YiS%�KVtu���j���t(����&	�B��$�oj���-����o"w�(���U���F�'���U"4�؍EF��_X�Qّ�����G?�b�Ԧ����e>Pe>�C��+�.d�	���8HI�#��gB4����ߙ:��2A�!#��4  �ma��'�b�-� ��%́��Ly�UI��*Y.k%��.�E �js�Ts�Y��x�hX���U� ��fn�"UZ$��[ʡ�FDP"$A���A륑ܥ`�U#"�U����(�4�D�iMش���h�s��nX5( ?Q"!���d�ykԘf��"ڗ4I֛Za�S��'؀�r�C0zsQ:vY0@u�$5�ly�g�5��
7��d2;H"�H����:�d��̌��i[���f�]� 3� ��)�v	��?f���KJ�I�1W�� r�ր�x���yR�aD]@�8�����@��d4څ�/�%*��Hk���]��J
��(�������I��D��^�]����|,�%ѹ�A �0H�D�@�@��	wp����sϣv���`0���r�%:�M��(�I�j�E�oD$ bp�i�_Aw  �  url��O/l��R"e�Dle��HA��z����Xh�v�Տ/mu:���h�S!���@e��x��%��`0��U	�Y��l�ț�R �a�rN�c��#0��fKJ@�b��qP�^�Z�TK�
� p�[����m��m�م�{�f3�r����V����)�����