BZh91AY&SY�q) �_�Py���������`�z�k��� ����vt�{h$��dS�4�mOSM�SL�1A��F�$�M4M4     s F	�0M`�L$�D*z��      jQ�d�I���0�� �2i�$H=&�S���Q�@ 4���ɂ���"@�
����B�?����PV $�)��b�O� �b
����J�@`�,ζt������K��9��]�����fffe����ffehH{� �~��ɤN
��`gwuZ���1^�B��LT�R)�Q
�[
1iRH.�� :�-��b��Z]T����8�~sOc�~�
��d�3e5�zWC3�&����6EK��[j�aUMQL-)Ჳ��P37��F1�	����+9��~dT�[�J+�<m��l�B��R�o�i�I,�ZxMW�e�nI!��7��R�e\8���c�z�-5��RZ�W
\�v(h ��E�KI!ٱb4�2��8��Iu��m����u1k��� �6�-���G�rg�ǚ�џn����Ơ7���OL��'{����-40n)]@Y{0$8�zᥕ��S������%lHK��ZS�y�L��*Kָ��`�l��U�)�vW}t��� ȇ��D;0է(I���;��� �*\MBJ��uYF��N�j���Z_,Yi�K�X�xb5���tX-єP@$ ꎘ�Z�M��'4�H���.��,��vWN/eMn�1��Ѵ H=��b����	���k]d��p/�Tx�{�s���V]��ëWTU�r�&ޝHnW�r���G�9��}-QʶAeڄq.�l��09l�wM�.X�˕�Pu�F�|DD޸��t'�Ǫ��E��k�[�;;v	q�ۑnf���#8q��<�"��+7MW](�P�2]`WR�yNnƋ�{�F�=��QWyVhNG��I�h�w%iO�Lt�$-mzuFS�[*�-�~�V1M�v��2�E����[kW��`QA�4hԊ2�[) �j�������LL�����\�WDD�U4��j�}��7�e��0Ŭ�V�&�!���b���G���ºtz�i����������8��ѷȋ@"�I�F������R��n�߾���O���kͮ�)�عr�$�ɻ�/b�RӗhXp��!�@:�� W��d�I#�!�Mf|o����6P=��$�D��#� ��uL�rf��%��@h=� �(��ё%��m0��%	A�и��/9����U!ɜ���tof��w�� h���B��H�-f�X��g��P��vk��
��0�� �"�ԩ@��(�a��7�4:]�XY��S�`�H��q��iU$�A!7@�n^FŇ_>����[5�F�|'�6k�X����@�G�b_��g�mJ=~�xnۅ� ��9 �4s>H맵���?c�Mw)�DV@�&g{rh$H�g��:�/֘��5����|�jU��H�0a��<��4�/�����!�D�3��� �0 ,p�И[�NF4H\�Z�I#�7*�20h[	%߮ (F���rLl��t6L͉%S���,rK	��Ж;�FʪVImJ�X"J�Йf��DYy�xJ�g��
	1����Ո����ΒG.�h_wv�P!C�^�n�z`�B�Z�5��|�m�%�sO��8�d �P���ï�8$��I"g��x��|O�ĺ.��2�#R*�m�@�rr�3�3����a��^�J����}�}���C��%@te��""	�܅r	�O]��H�%����HYuv�Я]k���IRV�ADW�uz�P���k& .)�1��bEL��$���9�˖ [$��
K�����?sz���F��Ʊ���OEn`İ���.�p�!~�R