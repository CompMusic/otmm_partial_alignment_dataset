BZh91AY&SY� s/ �_�Px��g������`_{���;�z  w_��r��}�	�dO<���4�L���� � I h�     50�S!�	�	��4ѓM4j"	)�d�4�Қ4�Ơ���hh�L���1G��C �&�ɉ�!��E#L��&��d�C � z��4=M4�e �|s�� �^
�Y �\I{��EY$�RH2����݂HM�	�CR�J �*�YO[��oQ����x��>��]��݋���̻��������]����K�����w�aҼ��F��vf�ҫ2��u�\+vmEo$�z�r��+Ux\^,a
b�0��$ǻ�bT�R�DL �&����D畨�mQ5�[8�8L[������-1��)_ DN��7%%�����S$2}T׌>�j7mqۓ[T����K�FE&A��*�x���i$4��>}�6Q�����bl�p�#2qAY�%%B@t�Ƀ�26dhR���s&��SI瀼�Q���ix�>r�75���1$�A��Sd��a��J����,�}2	i
7*â!���*,�iV��
�����d�%��C��;��Up�t�^�ScĂ��_JH1J����ݛ1�0l�D��/��*D��F
�C��,��B���d'�I�l��(,�O"���M�h(˲n�b\���oZD�A�p�t�K�V�����%Y`t��Q�Hu	�?
庸r�$�����!��e�A0�����o{<�8���BIɀ6��jTS�^GT�O r�B��ӎ�,iQF��E"���s=m�
����+ki�ۡIlU9|�Gh6�i�7,��]�hE�\V^g4IW������J��^=�"�H�½N��.�$��#�:&����{����q8q�w��w1p���.<�$!����`�|�sb��Q�Ȗ����*4��Ic�Mkm�t�TE몪hNo��<E1�G�Vi�^C9�$.��}�G����PS���]�p�]FVE������r5�mE�꣣v�h`,A���dX��*�ݖa˖f��+j�E�b��DI��cfws�e�a���f��Ie�h�ћ���O!e/���R����۸@u|(�ǣ��UZ��ꍝ��М
V7����g�o��.�uZ�rI#�>�N��T�����ag%!�|��2��U9HR�uƆ�>{��sK��O��S.��A���x����};XU<��殃7tA��Q)&�C��d�q31����n�q�t��ػ��^BG%iJةD�5�:8�a�q��$�.����`h�
H(�:�QDEb�2o`9�Ps��FU����8"���r��� .D'fL!; �2)��S�G}=ɀ�d�5�ԈU9A�$��H"�3]��}kͅh�D���!BK'�9g֬�b���J���=��|�$e�;�e�vG!"��^��_�!��mI"�ɀ&=j��A�t�ߎ�����9�-�M<"���*���&n�aZH咦��*��v�1	j��[���q�1�� [�a%�BZ͵���K"$��,x*�Y$=u0C��K�'��:`(�P�L���P L���X�~D��TU�y�P��������Cs��)��ÿ�� sl�z��4�5� pj ��^���T�*��΢��Vu�pDd��y�+���鸴<�N�S���tM��o����(L��쒌��" �~�������3BQdI���uᰶ��M���IU�*Xi�q�!����b`��1�,�)$n(O)3IP�` �l��+�G�اVYA�}!�38x��1,�Y9�G�]��BB ̼