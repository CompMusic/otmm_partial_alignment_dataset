BZh91AY&SYgJ� �߀Px���g������`	�{q���`� �0���"�)��0F�4��444 �)F�M2hh�4d���`F�b0L�`�I �T����  �� 4�ѓ �`A��2`�D��#A�"zOS�jf���=�4�1L�x�R!P��@��^d�EYY P�q��h��Ȁ�Ă �A =T��@��Ow����&#�2�D;�fe�ݭ�7wy�����wwmwy����P�~��G�K���Au�u�xX�BK�1ḽo/*Ih��S :� ӥ9��@�-��R���4�ul�gL�w1�;��B�,<�]U��0�D��aR=tY�,4�i�at�u�G�S�M�+�A2F�H������Y����9J%n�y���~���CǦ��P�&$�Q��J�JEi [A�+J��W$�i���y���׶���tkʚ�ywed᪥S���;��R0ӭ\\��b����[�Exюa���.�;3��>CA"��Ӳ�J�"ڮ��� *���L8� �J���%�C,�G�2���E̸������Q��ha�q��|2�&b�^O�h���pIP=BW�z��@R�%
!#l������tf�P\K���ZBs�Ψl�~6:�*��e���Q��L"Y�(�U����Y<��OB�|�B��5�Ғ�ʽKD	�B<"�8��.�<M�	2���㠜�Ð@h,$Wjp�SUt�,\,%�9�����lF,�Y�;i��T�ɎX9);���H!�a�.���92�e�a�i44�R�2�d��Vl4�G���v��4��>Ԥ�Z��,,;k�����y݀덩P�m� 1V�ߓPʱi���U�Ğ^+�������^Y�O�e�<�H�s��z*�U��X˪^�f,,��ʊ�+�<U0�%�ĠCzЙ���0Q��b^�&��(͆���H���XZ\eլ��)E<L�!k&M���1� �{ϒNn�����
�!�n)e�w%��m����C�܆��Rż�Gq2u�*�4�^���̖�yQ�g�8� �}$�����-��|2�E��l%�\Dy�l��]u[�p"x5�N)⊥R%Tng#Z�'8�j������<����C̼�B����zUٽ]�ݝ�ru�K��|9�Ϥ�TE��U ��ޟ,;�D�W�̓f@�;^ܧΛ�Aƨ���UV�D�[J��J�����1/��`�R�6Q�f؎dxeDAPdRs��4��T`m��Bhf���+6xLkr�w
�j�mb��!��0�u���H��{EkK[&�A6�fr�غ��_<��O��I����kaJ71RĶ��t�u�I!��%z��f��!M/�%�
�g�ԫ�ٗ�9���/��<�
ѡ�I�2 pc�Q�.Չ�<õ[&�B�#�@8��̏. k�@�^�����x�~���62�F��zV~K�M�Cl	D �'�*cc1�������-<�X 9k7��6C2I���x�CK�
E���E��*���$�(��0�|( s��l���O��l�^�1pҚ@���D��*��Mp�kV�5*����V��D;���&����I��|��d�/N4?���i���A�Mn}ίZ��H~��^_z��p��iF�H����e�a���2��n<��[��M�r@Lx���|�%�U�Y�k�W 뒇^�UP� �� ��FG��ѮEJ�v.H�rU���i!,�̍#L���]0d`�H02d�=3t�n8`�ڬ�K3D�q�l�2��WeZ�t�2u�$ ɵa���OV(А�H<x�F  ��L��C�J��h]h9b9���x�᫾t$m��P�@ -�rLb��#r@�I L��U��
�.����E�*m6�8� )8����\Uk6m��p�mB�vs�
b�R��i�i TY� �%y=�W�3��5���uZZ� ��wY"aD����/��y�10@��$v��Ze� _��XY�f2�@h�6C��A�x���ڪ��Pc_�o�.�¤-@��q(6��H�
�UA�