BZh91AY&SY�Lg� �߀Py���������`�X��l� ��9�a���&L��������54ddC@1� H�       `�1 �&	�!��L����DT�j=M �     E)��S@!�� hA�"&��S�=)�zO)ꞧ����� zz�2ic��H�Z2@�>p�q�8X�  )U!��Q�*UFC$.>�!�Qp��-�ͬj����kٷtc��������fffe�����ffV�aaH�o�±��%��uCz1������iVW���u<JهKP���J,�u-0+�HUiDB���^[�{{��V�q`���Lu�[�IM��m�⛷�aiմ��P7��:9@���-�p@�	>r�$�����2*��𠹃���Iѭ��4hP��a��T�I"�"��X��j�f�CL������˜8��`6o��Ys�హoIη%(�p6��M���e�,R�S��1X�����Q��xc����;��&��t\�j��D2sw]���e�|�)Q�B��KFv9��tC���B�-2�"A�.�B��Ɯ���DM8���3P3]:���i
n5�,9i��8F��.E�=��֨Vô
B1�a�s���Y
�ʭnf
F<Ⱦ5�z&EÖ�A|P֬�������º8`��W*1X#HI(���q�p��6JV
4�be�tCݒzB1U �0R��F�&�8��6�=Eت^"/O��0��#�k�v	J4
zgQ�)���x܄sX2�'����m��پ�bף��8y	|Q��{�����1�e�X�c�h��ف%�� sv�ZZ"�stPp�1Vp@�`�"ۋ$�KA���!���fN�Q�z�!!�p��\�2�͙�Q�)����H���9��X�þC���6
�=��
	їk�qN�[��d���Exꨠ�C"r8;!�%:���r'2��fC����j�=:�.*q2RT���EdXc	*S,,̊�+VF��#4,,6��B�D�04б(J,2,�0�4LE5UV��	u�^I�,a��eDEV8XƬp��ü��CV:��+�f@�bLv'���wCG��l��-��B�T1v�Rx�4��-�O
� {&O�w����A�
�c�Hr��Y��(��*i�[�I#�7hG�s�뿔1�Y���ޗ� ��wi	$y(@�(�;���~5P_M�@�G�I�/�f}��e�{��XU2�z�rqۈ����������US-!�@v^��+`�u"�z��:�;�l�rsV(�]��z�6(A"XA�aDE�Ċ�.�pqs2��5��,�:w�iUI#�Ј`��?A���MmW�D[�@���l�bEd��$V!xsO�[R���_׶�($�;��o�8��::����JX-�������<z�vί�����źv7X�;-5�$�As &�O}��u����U�e�ѥO39��$���z��q��%��ұ�t�	�Sh,����pт��:�aR6��<	A��B	5�Ido�\��JE��#ӡ�rDC��C5&���Y`�w&�7��ʩ�{:�)$0�
�xq�	�܌�$ayBG^�KA	�~P�3�0ޑ�Z�5e���79�y�eF�izp�� �%-�#JIH����GMs<�+
ٴ�8�Qd�� aǉ0�7����D������G/�qC��&�B����*�I$��K
�C�3�^%ueJ'S�2�"�ǟV����0i$AY�0��X��z͌L��m4�ZFԒ;��ј YJ6 )^m�)��y�)bQ2�� ��e�I\�(@S���"�(Ho&3ˀ