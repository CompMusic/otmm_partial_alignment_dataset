BZh91AY&SY:�:� T_�@y���g�0����`?z�w�V� yFZ&�@$�4L��42���z� �&�К44� �     Sb�?ҧ�  �     	4��&���!�M4�LF�ѓ �`A��2`�D�'� 	=4�42  W���@�@$X�������{Cו�"O޾���BI�H��bIY\���b�x����em�`ҝkZ������̼9����������,����&��T�#}��j�"�H�sP�2��ĕ W�t5�o0$gk�s)�Zt�(��7�ҽ����F:��3WD�$X%�|�py[�|�l�&%�6�%U\��;9ߜ3��Ͻ�"K�O��SZ�̑�.�+2�Lx�6)��Ƀ�E���"�YF$��PR�a��$q�{���L���\�S1��&��p��#�e$�`"+��%�BFJ�%UF�3
Ѵ��蹚���@�gc�5�o0,���r?��7V:��V�Q�N�ҕ�f{��0�x+f ��6)�����R�ֹ�&3���+0��'Jj��
�r��wĐ�4�cx.9+�`�A����!j��eqZ���[n�d(ㅂ��U���?q4�2��ň7,���0 ��S��D���n�Ct� �A/+Ԫ��b�����zHpnP���K(L
ā�*J�J`#Y� �m����H�@M�I/̌�E�T�/,1e��ނ������[�Ġ$��,�"���B 6�"�-1�[���P8C'��֛�$N�J�S���Fw��l�P��p��,[p�a�"�<�u,�R·���v�ZN�
��t�X�v�rE��۷an�+����D"=݀�.���Q��8έ"�r�S�I ���Ɛ���4�$ �p'�¢��	
�S��Őʭ�w\u2��S�"�s�Ez������Q�؃y�֨�����Ԗ���%�Н�S�ܤ�,[�0�^%�J��VxRgg��QW�TR����E�|sk�͘�&��|L����l��#+D�-j�D�r�HV��*(���6�4�X&���8M�X(�8[$YL�E&<MQt�85������\�YAQ��Z��kh`bV���Q��c�K%�WG�]��?����.��
"��%M$愧.�U1�9hћK��(������t�\ʧgkG��k���9�@ l�����ݎ��������%�E�	Q�a9dָ ��v���Sz,�r��8��x&���*��������5���	m��#�G ��e���`ϩ��V2N�C" ��&� �X����4o����炇 ׻aq3'������w�;�R��I��lF*��c
zzBZ K�@^M:Z�_�Rt?&HI�Q˝�'��Q�����s��X����QL�v�Y3c't����}N�j�8̮�j�@�Q~�M�m��n�U�s����@���\K�5j/,QA5hZ_�r�f1�R�B7�U� ���y��Ē��gs�`�2p
=ZT	?K9웤�O4��㢵M:-N�`�eq@7�ƌ�%��#뚒�I9��՛֥ź�UiFљ��7�q� rGf�9N��B��\�0�ʍ�%��Q�v�k�Em�ёP���&�i�@����73�l5�ˣ�%��]y2����'����a�1��2ve�цQ������Z�Kq8�D�23f�b[r�4g@�z{�湣8	m�L暗 JR@�2A�b���)k.�c_g�h�$�e5�.���"�(HcB�