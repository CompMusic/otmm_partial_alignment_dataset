BZh91AY&SY
1  ]߀Py��g������`	�z�t��P tyNq:�u�cI )�ѕ=OM2�(�OSM=&��i��P1�@� ��	���dɓ#	�i�F& �&�"i5'��2i�� L� 4 �E�{ԣ���򞚇��A���FCCP�D�1S�S�<���ɡ22= �hh`�x�(pD�O��T��|���f��� `IC��J@��
D*��F0� !y$2��k�?oW����Tz����fffffffdDDFfffff���̬���GKE \��t���B��v����UL<�D���sBR��y=�E�4�=��8�XMQ�J���T�v0M�Dpp�9�uؘ4�9D�C�+b�<Dt�Bu�v_Y�r��3s��u�%-�]�U�)-�����a�{�;��֡ &�|��F''��w���qZc�%�D:��{���C�(|�(f	Ej"0��",*�^	&L&����NL�s�Q
z����H~�k�9�{[�Ym�7wB�f-eUj��A����5EV]��Z�ZV�5^��x��D��[	�zx����D3�iY�ǱWTa�w�{���z���h��uu�ӥ���
q�z �;2�H�F�%�B��
�QlE|h��[V�c����Uȸ^=,6g�2�hus���]�w�)�P;������ïD�P��ب�YO�"�p�qX�.�¯!����m)Q: A�����Q��(�(�iL:����U�h���wc��F�"�.�("Q�k�E6,u�Xr�[�Ď^l���l��u-n�,|�,��]����|��q�_�I���;rB��wu$�6A�� �%���EbI��I^�;	\�.Ð�@��ք*�n"�'9J����i��0'L_�ݠ�B������N�S��g#Cf,b�by�[T�����5�iH�ƽ�� �`��X���V�ZfR�%C`N�7�X�2�48�Y �����JT���I0MsB�4 !�0%j �M� ��5My�P�U��/������I]��,d�-��f����5������KyjL���b��@9'�g���2�;릜,ۧ�v��>�7/v��qww��Ꝑ���YX�
�37� ��8��c�",X���\;�������^�ڸ{���O����U$��r��0��*e��y�����Vf��j�Ʌ��AH�}F0D�)��x��R���)�)��AAD�#"��)�E!��-�
Ab�[�Zl�%�k�L�0qe2��T��x��=��p�_RL�i�l
1��<1O���yeTǮ�l#�����d!�!�г�z 1y%��XM����J��({]�Q����A�S����Iu&;El�N�Ǧ*�e��S�$V��<���I3 �
%����� �)]̇��;� ��b�&Y|�$P��K�he��\"_%�9A::h���
>�W��_>��D��"!�92�\Fʩ�?ΣX�\�q���இ��h�j3۬�.��O/�o�z	�2�����X*�H�,�Aa��&�B�zC`A΃F�n����S`�'��x��B���,(34`�w��8}��HH߇�!0m�2hræ5�-D��7k��М�-�kݭ�C����M1�����jv9G�g��t����MW�ö���[�ӛI!,����5*�L[r<򺥥Mv��e�$����aMN���ݕ͒����2�I��j"�� �K���
�N��HNnbq2�y!���9�����q��JQ��WKu0�QF��I+�Cq�h,Zk]��jq�,y�EU
���S!8���xsH1�[v]2~�<++sD�\�`:}d�&�r2�K�	.�U������&a�u����Il-椮|�t�%�z�i){4W�@�R��Й�]P+]G�iz&��i,�H�5�(T�ٓ3 �EčLPDIΏä��L`0�s���Vĭ��9�u�v�f2ϗ V����I6�[���V����(u�������� ��c%���$�_X��B�_53n�-P��������X��MnEf�A~
Dq�k�ʈa�ĭ �/d�.W	9�[<EܑN$�D@ 