BZh91AY&SYC��� v_�Py��g������`~��-  ���q�ˬBI&&J?S(��hd�C�Pi��D� Ѡ�   �	���dɓ#	�i�F& �&�BQ�i�@=F�P�  � "�j��jzM#F�� �   $&��H�&�4   dr@�]��E&��܂�B���+��d�q�"O�:�I&�w�� � V!]�ޓ��={yk�)9ϓo-�{�󵶪���.����33"��j=)�՛G�0d����U몠���P%�iԥ�����6i�Ul �CP�UPY�Wzb,���l����Fu󷯄�V�8��jd�e�vV(\�x0���m�to���N�Me�����E��<�D!������Ë��S���]!չ*A���{��SZ�Z��\)d1�' t��,�5 �Lc�͵uq�mUz���=z�'ߕ������p����c-���)��u�J���0�Eᗠa��j��F3x �Y��ŋ�I�j���m�%����NRۤ�i�(TJȋ7Ѭ��JJ2�ƋκKeb���*Zp��y6e�q��QElc�Nl �*"�A�'��'�IR���#8�h&D`�\�}q�T��~hA�fF0]��;�Y�_,���<�X�`��(0�[JcĴɆ��-�+.%�����p)$0ԫ�n'���`�Ep���7��p��Q���ɠ�����Ũ<����h��d2��m�A4�R4�S0e� N+���� �0���3�}���hnH��F��Mn���;`�:)��� �ɷg�Nf'n
X|Yf�M�cHz��� *S*+��_�WB�.T��.��Kht����#�q�-�H�3�W�5�rz�*�zq�J|x��#�r5�+��[v*:��=���;	�n�D#��;�`����F�%f�ͭ "GW�!GH�p�썡�2��Y����r�H�
�V��Ֆk'�C<��f%�V����T�J�Ć@d�B^�}��H���%Djy[�O< �$+�UA�#Bpm�i;�%�c)�	2�r�M��Z?IADT�
UVB����!l�RgR��!�Ha56�.y�c��L�-�M9�*"(�v\b��T�v\�N��j(5��g������2�~x�:�K�<z5��C������9�7Q9'��`|��e:�Cc3�����:���[����׭B
@%�q'����mdr��\��݄�6��83���73�t�����$���?xɦ/ 󵀵�]����?N�i�XD��d��ɶ��$�-��hޱ�	J:�H��n�@����W�)Q��&�ld��0`"
�e"��T��8`gtf��Xa�u����H��c�;wj`泬��fb"<�oS�a��, ��B��|���V�2BO���{�kG������l'k�CY�N��-�$LJ�k RTY���[�k��p���,�&�ƣ��+ឍ��]������y~ب� �U�&�6)M����u�r��k \�@����{��	ih �o�	�rSt�XX$<I��h��L�%W�,��9ꮧE[0(L9���L#v���bA.�E�I9�?wO+����+L���"�G@ޠ�'�0C�djN@�b[F4_����
 ��,tۏMʋϜ�۬ކb�pDٰ��lZ���u7Q�,�|��l�D�h�RXd��%�T�i2){`3���|^����0'�zr�ES\j���I�];��D�v����`�@�4�� `��L� %^�96b�	\��$�ܣ
ك�ߥ�z�k��rGD�5����]��BA^Zh