BZh91AY&SY�e ^߀Py��g������`^��o\8  0mގ���2 I)�����2`4#����M BJ� �� 414h� ���a2dɑ��4�# C �Q!)���P���C@ ��'�i�=C�d�!�1 @�� 4	��2e�P4�P(���Ru�rY+	k���D�]ꏾ!$���Z� �B�^�Gy��i�Ҝz�w����oU���˼�@�#6�jg�͡�:q��ӷJ����� K�өJ.!��Ø#`�љ5�	(�J$j���b�V�W��������Ɲ�k3��<��db8��b����Bg��ܸ[l��k����0�C$7)^�����/D��_D�BIfdv��?��\���z�H4j�yE���^�Zu.�˓�	:^�y� I�1�o���t�).�j��vs��H�B�%��y=��*�eyU☭���1#�z�U�f��2�2�[��a�7���i`ŋ�,�Bhn���1��)��0��hШ��ssy�e�%�4�4.�(�J��&)Q�h����K���F��g��f�mQJ�QJ��g(NȒ� K�=�	�`���F]��C,2��	y����Z|�rth9+�q1O��im#5��:�y�4�RrTk;n�-$��w��ZX��V���ɫ�M�=�&�F��ÓA����R��ƙ�)��ظ� �[�1�v���i�ށ��$#"���V�3V��OIvG�롈�<��W��eɷg��N�)a�e��0P�b��@
�ʊƶcAv�l.�%�;�p��Kh:Y��[
��q�-��g�<�O!Gl=8�JxX�I̔t�L���*67e���W�aО��Q�x��sx����d�., �*4qXw8q!yæ�܍��2���-=nkYq�-���74��K	;�c�pU�з�Q�n�����Q�ړ!+\�cM�I�{fx.���:a�7�E�UA�#Bs�]c~���2_�2�@��T�93B�-��3EL!J��UR��t)�Jf�T���Ul���,4�\�U��b��	E�E�[(��?�[3��E��Y���b�@	����_�τ\���������9�y�|�ܷ��#)�V����DB�JCj��{�@�'���r�4��[q����[�9,ʲf���w�[	�
�2K��0����Qf&m0�I�0L��؀��+K��:�[֥�{,��\��Vb��vKl����C*,0�s<��Y�B|�(���(Y�μ�*0���`��l ��P�*+AXM�A#�Ss+Yy��(��,�0�NO��[���+xҬw��t������NL	�_�9䓆���k��aE�C��k�k����5#{��&��s��+�ۋV�L�D�\=��5�-���p#0�@�؟���8Hm�.ٳ���`W�t��`�+�M��IEd����2/3��}c(6�/P�%�d�l��#6�f�@Jgn$B�C�"���X���,�*zꮧE\0P@�CR�A7kE /H�����߰YEk@j~��E!��d\^"/�(�h�aM��1Q+��Ʋ��-ބ�;���� ��dx闢��oY��3Z,6�t8� p<|����0�;1�l�拕%�
�b-� �������E2[��H%����H9깉�;�a��++�0��Kw
�����	{ӿ���'��Kh	h�*Wi���K�R:�B�����7�̝�1��:�s�	$l���.�p�!��