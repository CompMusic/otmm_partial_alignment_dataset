BZh91AY&SYY]� j_�Px���������`���]�}��4 407�}���^'gO[В)=�MM�Ѩ�i�bPz�4 ��M $�@h��  ��  &�)�S 	��b �MHBhhdQ�C   h���M�j?POPcH�A�i�=Cz	Dx�)���4�    *(���&���!d �vv�y�	I �!H}����I&��$��+�N�vS�-�wB0ۺ��x�/�w7t�v���swv�y���Nh3B�u���	�����g�����8���DA.�Bhhٶa#�5�š�W�b�j�/�Q���Y�3��w|��d�,	�Ŕ�N��l3��ё���:�$���/��%�qQ�GT1��->fj�Ƹ��TD��}L��f�hy[�n�.����CJ�SU3Y'^E��cثlYq6�42�i1:;�i!�^W�۝�/%5���g;=T_I�ԣc��Q�9�bc �%\R^+�g�bhJ�Q,s�Se3�v�e#�g��>]�Ŀ'"g[vʱu}ӗ.5��U��{�u@�!9�+�����֐a��$c@,��0�c`�$ ��a�]*6T��j��ɩ0:� �<�1^�^!\VvR`n�J�d5��4�B,��p�5���\�^X��e��x:�ܪ��M{��s1��i�Ц�w�,jKH�ˀ��� ����������|�QpI"d�����@V|*L��i+�-h�eV�ܑ���̬�Ї륩Xռ�t�S�OYGMs�Ig/+�� q&񶛜�B�^��`"�u�cQWNҡi�R�H���5�,�I�ɋh�6p(vuj����	.E��
�����@g�nݫ���r$;
�TQ�V�aS/C)i��rQI��#d0e�V����U�8�t��}�)��+	l���6�����[���Ь�T��p���>+�2Vre����L�O=K2�!�$bʚ
k�r1��p��G'[j��	�!�"�t4��RH�H������X����k5_�먊+���2B4'.��)�;<Eb���1D�mg��q% ,ɪ�ʪ�*�S,���*�J�E�#P�AHViV`)	���G!)�0ep�������l��MYk+��މ{Q?u�L�g/;`Cc6�J���;��X�P�=�����_ϳ-�_
g�Ր��eu�+�YL�ײ'u���MP�J��~��D�K�%��aYC��Q��wn�!|e�L/|��UШ��� �P���X�C�r�D�?}"B�b�1�x`f�z޸���k�~�TE��{A��iw��%LB�j���H�2���`�5�"ֽ)���Z�I����c�emB�H��dX(�P�E�3Ck0��܁�1�ƲL�%j�M/
~���;�e��AF�FL�|�2,߳$�j�$]���{�ٔ;IS�L"�G�y$����qՒXՂA
����@��#��uu�U�/�i�=%�K�6n��:�ImZ�HT�]a�3�[�C�*�!T�HL5jjyZƢK#�2�E���Ō��r�!pּ�2-�`L�� ���@��&�)�ѥ#"�����d4��M:_M�%(����$*�騑W�=�������S1&���5��1��3�,J���H		�`��g�t"�!o�ȃ����v����`{��Y�(:
�ړ/^��!��L�!�	�y�*97�3�@�:fs�E!×���bo�J��
��eZ%fL͑&6�$v�38�v_���	�f��X�,�Ҧc<)����!��`�.�.�_Cw�2`��A G��Q.c�����g$$���a2Fo�݁�G[	�A���!�G�l�]��YQe(�I
M�@sӑ�}����5�vc�����m_w$S�	�u��