BZh91AY&SY�:�  b߀Px��g������`�,x�h� =�q���Gp�$ѐ@5=F��)�M4Ɉ=@44�i��Ԟ��  �   sLL�4a0LM0	�C`F&�	�M�M�mF��  4�*"b'�=#�  � D�FM$�2���P4�4d�Z��_-h�j�(�D �	ո����A@�cP:,�`t�
����j���p�,r�����mƹJR��6˻��7y�9v�wv�����1��/�Y�z�������Q����%��y4BԨ�iI�4�HQz��l��hU*�TQi�Z�8�-�i80����U=�	��4h/��1�ǎy�I�V_Y�o�5]m�8���.���
K�8.�nc��M��&'[�˷'�E�TJ�����;�5m�>���|%�!�#!$��̏R��@�E��@��۝}S�HF1���Y�b���g>�����������Cw�q؇2K� "�5���2"���H��ٱ��n�E���!�1�m6�'�N�n�tb5��ϦAusd�G�Ht%�B����i͊�l�9GWAjВ�)5u�N�$'
2[�ń�n.��
kU��H�-"lP�_1"b�iZ�8dU�"8�1x
�v�Db�1�=m�:.��Is��A$nYIG��4�ٕ.�Rp�UAue�i�8����N��d�9�����UY��h,�^��;"&&B�i�6��2D�EWu0]�[n���B 4�3m���s���(�)�P�ݱ�6����A%��T����P�d<d܈Q��#�WBIČ��4C1�Uf��0-�bL�(U��N@��I�H��bV�\��e��q�h:�*��P��`�����5��Dm<^�D���fw�ŝ�hu�Y�z��V�)�M�f��(�PU-%HVwW�Կ�&���zY�aݝ9�i�"�+�hR�'WW��H$r%�^�Qk%Ҋ8�o���H��));W�:�k��NW�_
Ş	�5Ez�UHF���w����Y��y��k#����&n�֭m*�-� ,��$X
B�k)e��M�}eY0�S!��XIF(R"
-#��QA���a���Cd;���͜C/&��*��2IęM�ؽݏ����Su~��t*�;co�G�j��d�PT5��]ם����ѫ��A���Hu���10�E��PuRH\o�-��-�~�k%�*Cr���Ѷ�dA�(	A{��N�ի5��a#$@������+�@�[���A��(���Es�'l�9ے�Ҏ����֞
��dA���]�ܰ��W�����P�d+�ȭh����g�5^�yB��?*�C
I�
AV�Y���*�2,'s!�߁�c�Mi6Lb�ϛ���I�T��%) ��>��X�Ns
MelLM�K���-�Hg�q`\�B��
=�����n�����pd��n��P���c�(�Dn��W(�|����5`�w���AqAYi�(l��Z��<�B�4�HL6UU�:��!�Fa�,�PU�Eh�(��>�"wxN2��F'"m�k��Dʦ�K�*N8+�Q+�6r��:1��Gf�Xfv�A`��1�����UT$P��h�-칤�d�va��3+XOm�I�����nա4�>e�}8��Z����>|�QE��Wv����n�͋�� jQ��r'I
{ 7&R۹	pDHT��x���53PC�S�4�\H�?At�Zk����}����6I�g�D3��YQ�1ʩW�P�ӺBB�<�ظ���![9aP@+ٍՖS��ac		�§ I���RFO�]{	�B�M�@�%��0
9��&��P��H��2Q�-2'a��t/�B=5�C�\�#�;3����H�
gU@ 