BZh91AY&SY	�� �߀Py���g������`O�� �Zaф�=C	�xS����=OHz�z����~�mM� ��44I�  @� � �`�2��JzH���d���    � �`�2��H�AO)�Sz'�2��yL��4��hdz#����%�Qx���&w��	76�I�!_�?�yM$�h��c  ��,�����:���S�x{�Z����\��˻������ ةYګ����Λ
��-�i0�u��k1ڭ�3u��P��U��qGdU�.�����op�8��9ۻ{{�֤6�f"��$%�hKԲ�[���v>ধ�v�  ��4�Y�Y��_r���Kq�ٸ�6�L�f����"C��B����fxxj�!6?�\8�5�ȆC�=\4��Q��R�%�D2���	Jns�Jb-�b�adq�9ط��pÎ�(�-�˙d�;/9�]�Wv�w���hm�H���4Rg�	b����m%,�����*^�4�W�@�a41R�E�^7J6,��9 ��-�\i�wwf�!�F��;T��!��i�ʈsxA�f�	J�Ҷ�{�Qa\6h4�X6�^��eKK�ӎf8R��G҇��ܝ��\�Q �N�>Օ� ��C��DV=�b�QH��Xc�
�ѹ�.J��Qp3])[Y:�=@�Su�db�PUI���U�u��n[`�Ж Q�.�������fYp A�@3YIsʎ�5%M��td2��ɨ�QmQ	7��[��Jہ�C[���s^bmoe��F��;�		P:@!x�eq�AE�4�ڟ	�eM�����qE{��TQo��C^�e�Ʉ���̉�CK�'�T�SD�i&�Tp�$�hB�\E�!�T���E��D�Z�ҊR�y�ڄH�D����B��'6U֒�jc,|���˝񄌽��my�ٍ��b��v�c�����Q�D�&(gm<�E`��4�/��b;$�ѫW�5mW`޽jW��G���A������R6$"�z5��0�p�',cv0���!.C�p�EUw�p\�p�l�H�T�zw5��cZ�N��Ō�B�=Ar���3�Tv�ٶ=�+�A>J����h!��d�F������}P ��v	bҔ�
�(** �J()�&7B�U��'�C�A�\��!�s�B��fJ��d��e�f#
���x}A9W�ܙU�/��ed�H|����&mH�ȓ�nI���j�_��*|�R�v�He'�"�La(�y�v%tm�e�I�!5%��Usn�[e�1��	"C@�k^�d[���9̠���B<�Ū��/K"�i�d8��蠖,j5� ��]$�5P��{��º��
ɩ;�H-e9V�4�;��!�k} �4t�G���#��#!$C����:���Ƴ���y��c��.$�H�5>G�ޡ!v��w�F���P����~����]��$U��o�@�!��>fy��v׷�����mm!����A	 á�=�&����0*̯.���B=$�H3D_�ڥ������R��j��1��º�.HD���7g�b����ic-�ƽј���
����tY?�]��B@&�o 