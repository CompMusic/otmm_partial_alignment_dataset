BZh91AY&SY)G2� ߀Px��g������`��۳�� w�W&!J��DL�b=&�OSѥ6���?IQ�#C#�� I(�d�   �  D����Q�����@h4 jB&�Hh�CL�  OQ��12dф�14�&��F�h��4�4 �  �'��
��0Hp�T#���l�b��HD�jy��y!&� r&h(DI$Z������
��_'��*fg��ޫj��.�b"2r2�=��\��X&g���T��E�K��KHw�u�.��1/�Y���b���!]E��)4����Nö�H����e~l���*Ũ&� �dwjK*M�0���Ј�i3D$����"һ[�e������
L��ֱ�V��1�T.՝�*�
�,��p��lq˓T/�'�{�eH��6�ZL��i�P�۹����y�$����� p#�ˬq7<��-B5�v��)Uc���RD�D	sRT(\(���*�f�X.�*�4U�Jb%��,�Y�\Z8��y�H6�P��3�9�D0��$J�!eðf����HVR$t�YJ!�6�!G.)���f7w�8�	J%"�F��֍�XY0H�`mș��T�d��Rԭ��7�.��Z�4� s��cc����E��I&x؂@�KT���G2mY�SA^*9�G�UVq�i�"YRƣY���y��x�#aBY*�xF(d9G5GS��6^��NɷSۈI7ӈǺ������N�@���x�Q�Y�J����]�t5�`��'���ı�Y��K+�˙��꼤!�C���e�86z���z^<�r���>^�ʡOHv
m�StO8[Ć�Zvy�o�|^��C�ڳ#m�`��4�V:�B7y���/�#���U��ޜ�y _Xם���@�$2�a�*�m��0��77�No7�b��g�3pp��R�v�Y��xQJ?�:�1�Ki���Z���8E���Q����K�l�^{�.�����h�J)�!��z�1AE0�#�]�rdLT�������BcHX`f�S$�J`�EB�S��,��F�VoWDm��c5�T9$&bV��(�����J&�
7��OӺ��6��a1S'F�(�jet��Ť��B�2��;Q�HWwe����},�H�j:�B�`@�@���e�ݚ;������ρM��q!M��Q�`/������g��%�;��!�>A�fF�!\�r���'v��ϪL�Rʔ�'O-������d-���A�U�2d.e`�.�M�w9=e���� �@C����b���I��F�Cf�p��!~w���!���i�$��Ǎ^�h�>�F�+�$j��>D��K����2��Rb�+fWS:Վ�XL�I(cd��j�[�Cl�V):�Z,.f���sB�͢Bh��s�P��u�$/��k2.�j XH�f���&A�HK@�$m��B��@���i!{�&)�+MI�e���*�EW��HN��J˧B2k#G+r�$��|-� �݃(jFљ��~M�����H����e	!a��aŵ�B�(y��W����{�ӎ(��ۚ.�x3����	Ξ�H�^�j���La)@�i�j�D�Wb0䶐��88
����'ef�N*��A�*Ӊ*|ڄV��l��٥dju+��\�yp$�#g��a�8)f]Q�}#`�X� G.���"�(H��g 