BZh91AY&SY�1 h߀Px���g������`{�]�  `}�=z9eBH�F���I��=�������##@ �i��Q��M4h�   9�&& &#4���d�#�P��)���0&0L&i�
�O�j= �F@bh0� M4�h��A=5O����i�C@z@4zh� �~�$ �� ����{H_e"����J�߇��$�7�X� �U@��N��>�e�<^���o_3333333*���V]�ڭ�R�m�b�G��yM�8'��Vsv��!b��6��N��Gl�8m�Kc�����j����,�nm�[�}�P�Xbb����cl2��OAR�5ڵcf4�s���\��a]��Y5:/{Q�I��d$T���<й��j��U�ݦRt��;2�x�����%���gZ�@��pA%krB2a�������0r��
��i�P	��L�e��T��\�4D�0
�e�{�0.�Uz+�f�@D
�����5DG�%�����`��*,�H��l��n[�t�x%8W�p�Y�tQ�A�|p�\�C �8d�D��j� 	V%�GC�.
�p

�P��4j��kT�C��2�������P !8�N��B+K�p�x�J��{���nJ���Jɛ滀�)��*5Z/<
�]3�sg��V�R��o/�O"Ȥ���lJ�ս� Z��24쬕Q|�Z�����ji�k�$6iq]�;�t��~�����\y�R���pEK7��v7�7K��T0��s��ڸc�4�)�B�N�(�j��@VĥC����v�B����)^<�^s����뮊d�%�ޭ�E�����]���D5������/s���h���	��6c���ȥE����p��0{'h���Tq�~���g̋ٳ����Em5��.�*1�}O�:� �A/IUPBA�g��NXXu�2꽌h4�A�uy1N�l*�Ȉmey�*9�ܪ"��Wu��j�.qE�a��
U�M�a�u�vC*�IZ2mE�ٜb�,�P�a���k0��0Ї7��"���n�^/E�ݞCv�.[v3 �	�>�O�uJ:@�P��6Cj�귴 �
�f����g���#g�|�"	�F�w���͡���,)z"��i� �=+I�(�ZL�L;Ub��H^$e�B3޾C6< 7`�����/�s��Gz��qh7�����^��b���(���?�g����I�@���df�NTa)#rڸvc_3	�a�lI��B�b2�'"CHM9;�0s���Nq>P��`��AxҚB=�P����#$Y���L�s-�TX7�y��a�H-�2��s�!
^I+^kbT�� $Ki�z��є=�]��o��C2�8���"��cJFͮ�q�֯��"�f��§R�	퇎uzB)L	z�� ~|	mʵ�s]yoN��]�V�&pHG��z�hω��D4g"��b^��̧n����KK�&FM��ʭ��
%&HM�U(f~{x����mQ����"�SSeɖ�
s���d����B6�o��	���2h?^H� ����h�8uI{Y�*�7s�����Ṇ�.�y�e�"$���>S+�\��A�����uOMn��<�,QF�niY$�7x�7�mQ`��?���AMt�R�Fؑ�fOzs_�ԄP�؈n$�'z��^�İ$��t�[��B ������a��ؑ���mb`��N:�s	�h;�HG�ڕ�{4�F�#`$H��ٚ�G��R�V��n8�n3B�
ʡ7��Q��]��B@k�L�