BZh91AY&SY}f#� �߀Py���g������`?{su�r� ���C#Z�A$S(z�hhS���cԚ~�B0	�hi� I  @   `�1 �&	�!��L�����J�ʌC454=F����C�0L@0	�h�h`baB���LI��3Ц�d�A�y4�A��P�D, _ D����I����b�?[�?���@_�Z�̒��l��7���ۻ	K�,T��w7ky����wwwYr'4iD�~��x?(��7��*�&GT�]�ad-��i��Y��l��$֨����!x��x���F���K�
l6A]��m��3���fۓT:�[e�$8��ºd��>�s5���	Q;ƾ���%�ꢼ���\j{�nxk�i�-����/%��	h�TkF���^�bva �0̈́z����j�U�6�7�!R�`�;3��hk)����lD��%f�kWnq���C4`eB0:�D[P3#E��!�<b��vf�p��	��vSU_��wq�M������ȳ�)��.�r�t�EFb���~T,{9�GF�P^+�q1�j�=�`�d(,n鹽���N����w�p3�ȝ{h�8��AF<g&n2�T�U�^e��,��P��&dd9n�U��#y��&VI��~0I�-$p���<���`���X����;X�5��Hu��TG�V� ������݈����{G,Z��b:��߿.V;�4G �[;	)��c\'_��x����a���p��bף�������qDͻ�Uf�vL�KD1�vۑ��ue�xa�q�ɥ�k�Z�E�ň(�DO�э��o�Ćd�j���!!Ã֮v[���;r;�F��2z�Ŵ�Qc�w�X
�����h�t5J�2T�@�N�3	�rt��l>�DQ^����A�>��(��ef�u�1����]�k��su�����WJ���u&�k2���+v�f��jŋ%H�a%lYHЈ�l�-�.���p��*�lV"&*����M�g8&^f�����t��@�M�%�j�?���qu_^j[������~�m�2uca�fSߟ�J+q�|M��1����;�r���JPc��H���*�ݝa�������v'�*s���v��x2�]gv��u�5�;�'bf��	Â�`v���ڸ��t���W(}1X8%e$��BZ?��HB)2�]�{"3�<o��'E���B)�I��vT�!�\<՞������@�) ����b1g:@����: ��[�R�>���H["���&�z����ù�i����&&DA��$/��P���J[��Gz����~�d�@�^�B�8�O5�o��.�����_1����L5��^�D�Y"��1��U��x�赡# ha$0�+Z��,�y�O+.����<�gdhvt��o�'G��L�gB�)���nw�BjS"W��H����CI�$��`���w ����2�U�I�"I�@�~u0C$�Ĵ�I��0��si�E �u��bnE>o!T=�]f����΁�̽l�+���햣s�7�/����5�w�Y9�@L<9'S�U#�Q-T��Ռ1�0�Z��3A&ۇՌ�g��)�Ͷ-�l����,��*e7D�U&�f1ӧSA��4ڳ1mN�"��hN(Q���^�3��W߲I���x�aS�c�(u�7<І�S��eX1.*k�f$�y�6�#2>ƅX��}�O�]��
q�����"�(H>�� 