BZh91AY&SY��� a_�@y��g�0����`_{��Y�  Aܥ�Z���i	�<��zL ��	�h4�*)��4�b A�b 9�&L�0�&&��!�0# �I&���ш�@� �� Ѡ9�&L�0�&&��!�0# �"z�4��FSd����h  hh�HJ��! �(\���J�N=��<�ؤ�`$�k��	'A |)���DIUS��wt��^�o����~uW����͗w���9�ٙ��������B�t����ȝoZVe,�wv�V�Aa��8y��PhR's�[�ݽ@�ǦZ���d�@<�*��_�xc����-cT��u*�T�;�M�G�DH:��i2ܹ�)*�cE��~ ר����&*ℬ���S��?+ۂ֮UӝZ7c(��Q���e��l�� �&���F2�
����I�0���}+c����J�'|�)��=8�ҚR��ۢ���37��yE5��iu���kZ��mK���r+W�v)�ڨQ먷j��A��w'�9J�^5��p#%��Un`e��H(�,�c4�y��4�VWl������*R�Pr)��%�p�i��[��0@\��p`KPP��2��XV����(լ��J�r�ڍ��hvwb��J|X�x�7qT�*Է؋w�p� M����J�Õ�5�<�*�r��
�-���;]�8�D�@a�T3K(FK�bhi�W02�&��@M����3� ��j�CHu�)�p�n����¥�����
�XB+�qM��E���2��ޞ�(uD2w�8�{�"v*	�_2���ol@ThQ%�*,[6�p��Pd�q���{�!7�	*#֋5m�Ui!��i�:��y�1�/�-�^��\sJ�p�:s��˙
@�kv���/32$6�*��5�A1�ޘ�xFJܵ[@L�*6��z�P��	�:�TYeV��������.�C＊�!�66�8�4�o|]�E��@��Hң�q)��`}1}4'5�w��.]Ã�ч���3���i	��Ă	���F����|Ug?��u�Hn���eEUw[e�QX/����Z�j��+P�*(�;tf�&"�	�����D�KXN83$�!�$��'eۙt�v�S�燻�cū`���`e��ʖ<����t�_,����ɿ��>w⍼�>��*$�X��:���f�f��ҥo�F
��.��ȫ><�(܁,�T��#���jʡ�tM����@KZ����s �=��l�˃��V����idTx�_���T)_Y@�h;髛�̈́ � �T�����X��\SV��.[�nrj"����R�PY=����)�0K/�W�!���ڠ	|�IӷQz�&�W�yǦ�Ȍ��3;8H��)� %厢�C.��fG�<�b�!(h �Eq}�ԍ�%Y��3Í6��D-�)jn�	I�1��U���Y�k�����K���SL5�K�F��Buu�Y����fd	)@KR�F|�e	��V���7+3/K"�4	_R��3<<�ɉ%a����i(*��
��ҠI���dd铇�r���9�6��w�&CͲ�=(�.�eQ���gBJz�\m�[��f��Ӡn��k�����:���mP�,9�˞��F��d�=<	�ͣ��ދ2U���C2fh���G ��ƴ�1��6�GƘ�������)T�UGm�w ���Fj9n&qZ&����$�]��0��0r40�4>9�M����Z�%� ��S# �Ig��	R��^�7�Ű�9,��Hƾ�;C5G
 �lD]�rE8P����