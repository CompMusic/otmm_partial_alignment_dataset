BZh91AY&SY8�b� ߀Px��g������`	?,{]�p� �}�\��ݤ�h&�����4���d�C@1M "��a20  ���9�&L�0�&&��!�0# ��50���z!�2240CA�RB���=#COMF��@���  �&����S�M�CF�=@C	��=M�W`�X&�!@������$U�V5�i��qP4 {��́�ॖ�M���kٶ��M�t�9O3332��fffVb�f6ffd����̜�2�YB��Ř���z�bc��!㝈���ų��j�
"mլ�(/lE�Q���%�*��&F䗢e�qrʨK���|�igx=̿y31~G|��D����'\l��1p�H<�t��ka�L�
Kn�#F`ʷ��T����>U��<&zd����'�q/�{�������p�Rzey�/������� f�`�hcP�����0�٭��ӔQa]�.�)49܍0�6x҃{�1H��E&f�3&c�����>�DF��sc�/+��&�E���L�O+{!]l��xav�3��!���e���AW�Q�sAX,� )8놧LH��H�(�'XRV�.ք����:`-���:�gl���RX��.E����ǽ�\bL9 �g��ź��$��2�u�� m�"IaPIJ�p:�%B*
�r���D�����"��m�hV.�d} s�V��-A8��l��=��*�j��v��l[�i�.C4)2��s�g!�=��dh�<R�kf�����N�k����K��u�"�e���<���R020!���ho���(�s�J9�@l뺯0-�2�6@bd��$�-������K�UpF�֨bٮm%�KU�{Y�%r�5lM�w��P#)\�E��}b�/䜷y"w�k����)B^(�d�Ӡ�4x*%��T�,��n�Zg�"0ݱ��9�!{��Tޢ"#0��ī�ffW���ｙ��V%���ZQ�� �v��F�f|�%�,`R@�u2h�"����87�rv��S�οzXt�^�+u��u��J*a^�p��e��nU����\���K�:����{ﾾ㾢(�eUP�(�O/�Tb}G���s��eYYS��}N�*��� {�\�X���-
���
S���KH�B�)F�2��Z6�5X����(�����Y86�H"��#�"ę7QQ��BM]���դn�����u�(�ɣHn��Ν� 85�:Ⱥ�{�Z]2����Ҡ}���ۺ��	^��N4�\�1>�W����'��ҁ���/�=��]	�嚏��T�Z�ɑ3��{ ��9@��2� �,��(�h4wn��s�ux��f4�I_��Ij�x`o�u�K�nI%�^�9ud���U��AUI5	"�B�hY�?7*Rvhee.Lq)|Q�$��|�CR��I*��o{>��Z���MX��
-!JB�� �KB��cHЃJ)F'Za��Fe��C8^�~4�6N�F�b-�_X��"5n�c����������{t��R�6�5W�̤Ꮟ���s�ц �pE����m��i�)@v$����|E5$Q��Z�I)@��2�F�ƗV�I���$�, 6�CW�����t���0VbZ�H	[b��k�MK�aJHnȡ�6C9U�0=�r�:�B �N�D�0_.N�ZQA���ý�d�[��A M7����b����a�/huL�X�
K��n&����N�[k+&�yssL:�]L��4�9�Yo6CzÁ�q�0#�r9V�_��>?�z�U��t�%�s(�bA�%�"̚cn����s�l����P����=w+���i�c�I=��Ut$�Z�
��W����i�X9��k��Mb�FV΋C���M����0 <��\���H�Wl��;��'@ X����t��=�,�G�+��:��09��������)���`