BZh91AY&SY��W$ �߀Px���g������`���6���|�@<�yU���imS	"&�jzh��'�=2jjЌ@�4�H� �   d  1"��hP�  �  %=$D��@  �   F��Q�<(4     	!��)�Sѩ�I� bh��d[$V�;/*$��,P
 #i�M)��P(8 �j!����  � .�'c�X���̎��$?7OW]��ukZϭ��wU�wu�wvn�33/32������P��f�����/��'�	B�c٭��Q]�V��^��j��&�.(u�%�m�-��n2��0��ku��y�?��"�BY2{5_L��3"$Udl�fTW5�h����rх2[��2ASqċ'��nG�eW5TJ��"�nϛY��Owb��g�͞�Ei+�f�(0v�v� %d�H�G�k`	2d�6�.;�r(2��J9jζ�-�jыT�ĥ�E`�4�3-J�I�",������X[�%0Q��#U���a�=�;lsmDJN����Y	��`8P����MU@2t�8`R�	<�rS"�*àga�u�#�C��k_2F	!]e]O�Yx.� ��'�  ��!l�Q�4Z(����X�Lم� ���f�:��
�"��D"��0%�G828��l�k�a1F��ݻL���B�qPF2)"��#d������`@gRN�
��x[���"8t�8\3��.�G��b2Y�`��-"cj��ґը��hM��fi���i����!H�ax�8���0�qa�K�CSX³z&7���2Ls�%ƍT��Yc�\ʑ�r�KJlaS��P��v���ST�� oWQQn��0��jE���p�ذ�{��&��[�� D��i�p]Ox&���`.��/�mu(�eu��4���Fr�y� 3n�N�x�SC�t��$v�u@@t-1�]��B{7H,g���5=��*�[��ZR��ܺ<NM�lm�m��4	8��˽����J�FM�H�J{���GD�b�q��	$��0�8��	�P�2�H� ��Eݠ���4T�e�	%"T�D�hUk[%储�#c(̆�ˆ�Ķ�U�[�����e٣"���W �6Z������u�-�7�ۏr��q�9w��=c=mӨ5�F�/���/�(�TP6)�Q<{�%����ק�	w*vY^��76�K�|��K�S�kHCh_" p�'fq�da��;`��5C��V�/1�O�;j�]K�n.zs�|�O��ʢ-D���\זw�M���B�V�Ї�~�&��z�XO~Ed�[Bf]Һ���CTo�j(-!B�-
����2�pv� 4�fj��1��*�˸�\4�X��ƄC@�\�j�rMlVw�ֻ �I�5ø�Y���B��+�K����4��S�K\ύ9��bd@���Y��#T�k?�����t��DU4hH���P�8U�8Ș�J���+Q��raY�%@X�c־y���Kѝ����N|B��$�����w����`�(��$�Z�09�&	HK��f4�0	a0�	b�YkWQafR8�� K��ũ�(,`�	fLjd��F+&��(k3�'�F�d.��A��c�BJ�q��q���,�RfGv����qxY��s�/�:��TZЂ�|�ė�\AH#�p����n�o ��m6�:��
N��C���滲�V.*�X�֨P ��U@	Q���D�'�������r�KK������NJ���*i��$[�ѱ����M�@�	f�h<t-;�,޶b^�-�D�%#�ٙ6�#�R�[Q�|c��؟�4�0Q,���w$S�	�r@