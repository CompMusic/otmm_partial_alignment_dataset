BZh91AY&SY�~�� �߀Py���������`�����}�x  ������N��;�Q5'�f���2i�4��dad4��� I$�1  M�  jzd��i�Ph�   �  ���&MFM�h @ �D�je=$��5�zM�e4h 4� �I�LAiOi�'�z�  i��h�h#=��%��f���F�	O��.(
� �A����E }� �^L��M�J��0k� ����c���_Zf�r����^fffe�����ffV�av�"W��3%�r�5���ک����H�uW��)���6R�-�"�l�L �T�i�	�"$L��i�|�m�>6b�p��52zczTͨfq��
X�d�Z�Sp��q��S�-1ک�b�`bn<��r 	UWH�R��]�3Y
�#�/��kF0a��\Mdݤ`�BS+B4���/�kt�`��{����4�Vјln����+�*�J-@��(���PpV�PMfS�	�y�X�D�%��Z�"	XlK��ȱ���,
rF5��n)i�]��E�Ȧ����V���e,�}	i
6�8�(UH�TɎƌ<�tI*B˺+�����F'�I�|��v5����t��`^�60�lO�U� f~�Dڇ4C!:�]���Ϊ&��5��X����U��x��D��B���dU^I'7�6�B��@r[Y ��
���9D �P��z���ô@-�8�OMֺ���Q�zX륔uBQ�8E���yT(�I��!|����m�)uA��3�ne���`X9l���D*��<c�@*�Vf�a<�WHR5�㭋TU��E"������D���vI��ǥ�J[wq��!��T�0[c������#�˼扂��q�3Y:�B�/�a$T���t~-ʸ5щF��]f{���b �OR�F3 �=t�qˋO9cέ��v/�}S�]�&B���eo.ui���i��Y�g����QWqUR �9��x
N��5��iO&�&���$��U�WѢg&�L���t���p�]FVb�JJ���j��3��b�G�h`,A���dX��*��A� 10I�Y`�C*& ��\m�:�j�g�P����������,}�I��sO�W;iŖ�QE.�t�k�ƥ�,ʼ�,�
,_Vؾ5؛���(W4�&��w�jәg�IhZ��G��UVI9��7���{����%�yu��!�"�Pz�����!$�p@�5�����2�|h��3
	-i����M������K�p�Σ�&*�z@��}��� A��,����~b�Y�)�&4Q��K{�(�Z��V��V�$gs�f����ʌ%$y��x��&�|ښ�AIX�DV*���x$Ts��1Y��S�`�t^��΂-UM�)!)�$�y��#�y��y�k�>��4��H'0�;$��؄WϚgⶥ��pݷ($O.�ARh���\��e�M킍B����$c�`������jkz�C���pf}Aݔk]����^��$�Cs 6B��$ݸ�=9����c>��vg����ي����	N�"����j������4*�4]%���3�z�i��!��(H�Ē��h$\���)�UC��:DR�ES�F��oK����-�T���,���S2�
@�Ֆ�ŝ�	��e�j>�M�0B��_� �6��2Gz��!����?�4�/F����* ��41��.h��G0�I>���+���W�t]��1E��*�Y���*K����<�[f��\�i��^ƞ�c1�貥�R��ںn���[qJ.鞗�n���,\��Ƿ�}z�r�v�D���Q_Ǎ��^��lb`�O�H�S؎���$�¥7M�, ��6 )V�3Ŵ~�J���F{cA���_ n��]��BC�6�