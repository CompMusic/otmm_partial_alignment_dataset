BZh91AY&SY��� i_�Px���g������`������ 7���J*�$D T��h�چ�@�H4�zji�i�H�L� �   "�S�=L��� A���hha&�)�	�4Ɉ2i�@ 2i49�&& &#4���d�#�ЍC�0�15O)��CM�h���M)����� & 
����:�M$U���!T=���tH� O%lhB� *�M�^}�{;w7^���qu�V�����fefffc�Th�B����,u���!x����T��b��u���C��^��97yM�tĚd5���z{��p�jXH���?m�9JG�{��a�4�J ��\�M:f�y�r��&�]�<�ܒ@/S)�$X��q�j�t��8C��(=�ҵ�D�I!Y��v�=~��Ը$!���]>[��}R���%ˣ,tL(��)�c�Y(!�)D۔͓f�6���1n[u�tf��gj� ���г]��򊭉V�:g���X�`�PwFզ�jt�	���������sL�3x9�$�7m�p���vYP9MB��g
�UA�F�(q��Q�gv�yͰv�b�����,��uW��pˀ���i `A�`���7��KR:2$],�۩��ڗ8�i�k�P&��Ur�D(`��dsC�Ǉ8�ف�ꥄ�2�ZĔ��0L
`��A
��R��[a�¤F�*��
�JO&�sK}E���4J��P��֠wL~L�Iӆ)�F�TYr����*�Hp�u2�R2P�����X���Rf�*k2�0�A=e��YE���(W�i��O+ � @cDt;�n��VƊ���Iҗ�5���mU��@�	=&��,�ِ��J�<�E������P4qs�Y�QW���! �;��Ϫ�yw_vl6�A��S�y)��w�1QLIY�lY8�PS4�͵!P[b�]ZE7���)7l�ӋQ����K5h�h�Z(�t��g3��E0k7r�`&��j��|����T:��im$@u$��U��d���%"�Lk�,�V�"�5CU+�����:�Z:���T�$HC7b��>y�_?��x$Z��$�Ѐ����p�ZalCJi�08���ZB4�_ь�8����^��QpK�ަO���bd<�s��T��������õ6�׷���J��N�&�y榠�Ąg<24�#s��4Kg+���m�s�F)AdD��4d�B�����{�Yk'8���I�ՙ�#�4�v�!Ӵ=��\.L�)�D���.�Fb�j	���;a$#�q���_�R?�񞆙 �"Z�KS���.�6)��E-]�����-�1��c�)�rEs*+.�lz�)F�:(Y$#0h`��оy�.��Z��m�`@Y��h@�lHG���^@4i�8�DCF�W��`��C���h�#"��"���ld^ڕ�F$,N�e ���LE�^	�jc�"����`�T��0L�V
r�SN�fwqD�2m\vp��Ԍ��Q4�ؑ�c$��wRw���+�:
˝��`�n�6�˜�$o�B��Z^�/��1�c����HD�o�MwW�u��ŝm6��:�ƨ�'[��1ճ��i�P��	K1V�P��jB(WLD7��
A�r� �r��gAC$!�!�x	@�H�g�W�$�#��D�	t���HGn�*��Z�0����D��`9R���֬�,�c_�3�z���4�b*���H�
�:#�