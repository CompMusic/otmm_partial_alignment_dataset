BZh91AY&SY�x �_�Px��g������`	�{q�����  ��Ie�Md�BE	�h��aSf��SM��M#�A�4i�f�i���%G�4 �h�  sLL�4a0LM0	�C`F&�$�S��� 4    @sLL�4a0LM0	�C`F"@����M�OFє�j�0b=54q�� ��@�$"��@?��d��Y@T?O�V��ԁ�����������
���}����.��Rs����wf��ڭ;���y���������������8�mT8p�؄	?^���+�*&�ǆ�\���(��L���SV�Qw)۝d�� �]a*E�k]rNS��D�ɩ����73^���V
ԇ-&�R�_N�<��a�����L1�XT�6�9H�4����
j�1R�I2M�\$�Z���I����Ľ��45�	��k-U|*�F]bp� �\����ק�@0cp}�[_7���j�n�D��w���$�\O���:ִ�o]kfݚ[x&Sw{sZ�L��WwNml���L� t�z|����P�T�</zA^!ow��Z�M�!��8t���u��x�,��@ps��wvs9�nl�[���k2b����H��Y�Bi'MJ�gs1����c d�Xpi�.`b��c �"�*_��O/�u�7�i�yB9�~J􈲜 �֏d�B$
�kxäD�O%�%��R@�`]���{�iR-���4&9�L}�mR_E�Uu��%;��o��#P��>XW[d�j4&��Q�s��;r9�T���u的�[�>Q��w�Lk�����4q�Z<��tskt�+)��*��y<N^O^�Nc)m̝�l�8(���+c)�?z������rdA�E7��"�*��9h��sa��ɩ���S˴&�E�*ЮZ.� m�I�7��[��ݔ�w�<��4�����G�v�a^��7&�uB�m1��au�e+�
��쌾UMw�����:L{7�ݦU���$6[eN6��{ۢ#�-k�mu�tDa �XM��/*9X�#��Bx ,=�;?������_�*�ĩyY�e�H(�\�h���C��N;n�v��"Gn��zŭEg;Ψ��N`��A̎��!�R�U�ͬɡ��aڣ�?� �knb�1�		-�+@����C�+x��]��͛Hv/����M��&1n5��V_̶�X�j[PYYUm��R�/6�0rҫ"�X�<Z/9�L
����g4riZ�b�}0�(��%)��e̯8Y�pj0D2��fvZ�p��G�E,μ�a$&�6�j�Bڡ��<�������%�G�U���T���iqRx�8yP���Y+2����l�󉅄���p��ʛ9�Ub Ϯa�Z��)e�/S���/2@����`x(I�w-��j3�R��/�&�Ix��d �U�=���%�~Ɉ�V\԰]�tu��ʈ�"�cH؃��z_Y&Ɣ`A��\��{��]�N�̍t�jx�@���mn�{�ra).ϧ�_nYG��shTb,��b�F*�TUb1!�`m�S܁����ٖd���g���9�1( �B�J�:[�*�!z��̸��
��B� }�Eo;��K�(_���=��eɐ4�%�bA��Gm9ݻ���:�z�Ӷ����4H�E7û�հ�Mk6rg�q�7�P{4B����س�`Ť �yG_�P�ZG���,�k~����e�@@��x�>=�ޓF&����A�
,��@j��h�.i��� ���i��H��@�T�bH!m�H(�t�M�G�0imT������t�)�2̧"�i�L��z�c�V��=x#P�;q�T�Ӆ愐a�˟+�J���$��_;K���?hGT>�&#R��ۖI$ �ĸZ7�Fb �
g���x\[�,,��8�'�l���$�I�&ߎ��l1:��ق��Wi���.TR�R��e�P�*`J"�>e�$@O�� ߖ%p���e�@*� D*L��h"۽]�,@d�˴4�X`�0=_+�lɌ� y.��$=�3������-u�5��c8F<��"��[����H�
 u�� 