BZh91AY&SY6n1� K_�Py��g������`�{w����  p7yW5dhY��A T�M'�4�B4�hF�4��h"��       53S!)�)�j�@� ���̓L�=&�    �	���dɓ#	�i�F& �P&#Q�Sjf��M2h hz�i}(-������`�Z��"-(��\���D@-D�Js�xM$y�}.d�T9�L��8�8.��ٶTKf��s�^fb�]��M��̻���k�̽@Х_��iK�\��i(ޅ��UE!'k�D�%&Rh�Al5+�p1׶�B E��(�-�
�TRJ�Dȩ`����G�$L�A�tg&	��l�4����30U�;ڊw�X��R�T2�(F��!{�Z�m�{lh���e�M��"ЊֹWy�'�q)�^�#u�d��~�-�E�Y�� �[i�Dͱ%f�P HR)z�Ą&L3w7ѓ6�3�D����/�|���R����:�� 1 ʸ`�
)�e`�Zr�G��%�A�μT"��{�.N���m�X8Upl�"$�{�y���bX�FQUa��u�wӀ𠪧��/Z��m�RG*{���VҀp�A����@b�aP��		f���P�xÉ�"�g1��	zh�ÏY�/K.���;�]ِa
�u�|�@ǝ�
|D��j�u���G˾�-��\�~܊��$m`���s�7CY���h�D��S��܅���*L��Œ�o3�oK�
W`[A�M�ƈS��|jʅ�$�4�~R�q�;�A�aظ'�1g9�'7t[�f,�dZF�l¼����]�R��=��$��d͚��j)F�j�:��9jf/cU�fu`pJ�Q%0�����9uw��h�,I2b��$�@��C��(`u�*����r�eBX��:̡���{��k)���*:ŋ|���c�.lr[Y���T�8y��א33�䎒���+��s_��v�� B6"�dS��t^�k&�Gl��cԛ��j��/9;�;�%�2^��lI+�$1z�s�����j��"9�g�0�X�ziʃ<]��iV�tJ"��Պ	!����GE�/��LVU'y*�_�՚
J�L2�DbکT����R���|���U�/f�k��k$�"�)�H)r�͐��,��K����f���I���i� ͇��j�H@"	�\��\kď�&��ew��;�6���!�����n��]�U)�T7��Qwc�3��47��dy�+�����(����X5ų���Q�[���齪U"v�Hbp9���*���pú�-kv`e�\�B��.l]�oڙA���O)�����Ά�c^\��!DHWht�Y��u-��^�]sUPQ��9�ja�~�B,�{f�ڀ�@0ZP*# �`��*�( �3����!�\�Q\S>*�+Jw�9�a(Dt�2�=��W��ͪg�Vzf��x/�)�Ne�1�X�Մ����{�q�Db�v� Z,�P�M!�lG�;��������4>D|*Hͺup�"j3"XD����i�֭s��k4!X0��k�/��1݌�^k|�<7hH��4aQd�>��L�c).$��;O#Y�r;����$"؆K���Z
i� ��d�w�X���Aaٺ�UJ��R�6d�qtd�rR��T�n�UiR#�ZqV��S2#�|�N�LY��u�w��8��DZ_ՠ��ÎA�(3Ө�8m��!qlԜ(���Z#Q��+�~΂��n\���+p^����Z�Ë�G���.Z�vG?T���'���̚�zm傱�@Σ+��^����.)���91�������U�HTߎq�L?ѐ���
��9B�S2#�d��1��(�QFMK���i�4�*~Xx�#���'f�C�.�p� l�c�