BZh91AY&SY{�j ߀Py��g������`�,y�p�  @}�N6%��a$�#B4)�0��&��A�2��M "�	� L    `LM&L�LM2100	55���P�=	�4 � Љ4��j42L�P�@ I$������h�S��5A� h��jz�K���.�&FQ�R�+���uV��I!�'�j�=��A��t3�,�@Qe�6����/�[l����:����������������̜����]W7�p�|]�F���pb�$+Ӭ�,������W�^1�ɫN  8D�C���b�UR�p��r��j;���wyv8q�ђ��á�WG�����^���o6�2BE7�q�g6�"�R�&]W*O�v��5�5@��(Q#�T�wT��X�n�*]��e���=�T�Un��2�=>���M�-�N(�&�r$4^�q�7P�]w�ᙰ���^�	qX�$:�	�L�v6��B���`��  q����([T�W��}���آ��c��a����������+���[R�tbJ���L�8$-�F��D2Ł�X�U r��q{�<;$�P8QD8�P�Jp��YT�
3�0����H%Ĳ�u>��(��p�l�-�`	�B��emH\Cm��E�A�RL��t"��EvE"g�JJ�3<�#N�d�+`|�\Y��Մ��8�1�y����� ��ʙU�i|�C�;6���2*���nh��'wf�V�^1l���}*긨���k��DX�a��rE�ӛE��]����Kp��E��h��`��:�D��1	S��H��S�{"�}�c^��a�k��Q�|K���B�P�����ݕ�E����%ݗ��9�b�9���jF5c
�OU\bS��YH!�i]��^&Y�G~�0���\R�|�#� r5ٗ^b8��Ox1�rۏɋ��EHB�'$Hb��#Ju��x��^g�)+`�  5T��O�]r�f���8ܐ<0C8�[�Ί����0�x�A� i�*((�+��fjY�������U���Y�i��l����I
��M��6�o�V�8/W;!�wE�* ��z~Z]u̯N2a ݹ�OQ����9�sF/6U�W��Vʥ������&)�RB�
���-�.�"�{fq���"kEZ�e�!��L�����b�(ɭ�Q�u����y��4���$�dM��缨����]এR�"����l��� �@�T87��&�3Q	L���ِ�EG^��&��;������*�?������4��ls�xՍ��߾�m�xU򨴞N��[@��נ���O�ܗ�W�M�U�T�(�R�ڃ�׽y[2)����f���b	ą������Tq;Ɂ�j��.eE�@�	`�,�2$Ԕ�A��K<2l.M��9�Xa���;F�`��Q
��P�v��M&:��rN��L�^�����2���̈4q�$� >Rs�[Z:|���SQ��ǖij;	��Co��H�g⑬�`�ڴ��T��g�cd 0�I56p�n�����;��;� �G��%�j�� {쿡F�3Z9*^���U,���9��t�FG&�\DT)Lk��� ~u0Lo�v%�I�f�#��w"��N8\7F�=(��_=D`�o�ωv7�en�s�Yz��u�Ø�Q���-����?q�e�j}~��GD�*M��C04Q�H���4�a��(��ǟ_��[��^k���]*�m�i�6˩�k�'����:��ĸ��/f�)c�-��ф����P�^�t[L�7���Y@[|�zY۪GEQ��~4�v�g��!:��p�C��p����)���P