BZh91AY&SY��2i �_�Px��g������`�1�[Ӡ�`���D�$�hjbh���OI�4h4i�3Ph�4h2��0	�& a4��R
 ���    	OI(���6��   h i��&�&	��0`��"�7��=5L�#�ѡ��z��Xw��� �D@��c��O�+� @8"0=��Z"�@��
@D(f���}?7������c���Wwwov�1�337wcwwgwq��f`�.���~���LI�tiJ���R骫�����*�Q��Ւ(ʅ� n0�yj'"�c
��#����׊Jb�+�\�A�Ù��%�)�TGP��ɢ�n�6�B�����6.E�\�䥂�Nk�Q�\��@�Y����ŋ��E�y���L��M��|�SJ?y����r�I�o;{{����:��7�W
v� #�D�ur�����Gn)&�I#�U��ZH�n٬��̯+w��[�{� ���h�+lm���i���\�do~����4��,���6�#Ȉ��,��ïn��$G��{y ��AYNj ����7�0��(�,x�rj��xo�д�����F�i������fZ�������c��)WSm�ǎ���wCPx�)�n�ua.Ƥ��p�0�⋽���f�!+��	h1��A��/�%���B<;��ʐ�bꝘY�8���Sl���[�d.J�"���}�'U_���W ��kWY=櫅��wrds ��bPC\�4aqU新��qkk��;-�b$R;4�߾e����������1]�ӄf#� ����c<����Wh��B�Z��ɡ���Q�U{Y�E�h��rb�.A#H��<F��"��0`�?�Iт\͊P�W�ثƖ��q� 1�
���f�8�6�5nd�,��M24�s�oju�lG2� n��Ҧ��#�q���|#�H�+��%QP��ݾ+S��=�d�E�^d{��U:@�s��1!56�"�55�D�����vG7�U˸�c��)iADTZ���Q��3p\%�"a���Ѯ��)C������#3�ߖ���(�s��xׂ�=E2������wd-���C�}0��=QnC��䨃giŃ�_H�tR{t�s�|ob�UhB�,�y�*wN�G��B��x����8H�L�Յ�FG`�+�u4d8��3B:���}B�����*Pԛ�Lw]j3T��_�.�Σ3#"#=Ч���ǽ�,H+�t�R�P�3φZ6=�`{�.�@T��J�mt��Z�D�AQ�ځf���4N^&!Ѽ�R��&&IA#�n|1m��pw&��PZ��BS��=I:V��&'ـ�q�؏U93T6�(Gi7����ĕ׆��N��I��rv%����hB˙���\�?,�|�͒����{�y��x�*������!-�,-d ��DG�s6`@^����Q!8I}�ӕ���Qr)PWa�r�j��0]`���^�PT��%3�)|�Q��ͯYyb#�k��3�u�4�"��-@��?�������X��x�՘��GPc�@�*J�L�7kf� 97�Mh����vo#����jp�Pn����fh#N���3�g陣��U٥��}ѵ��]�b�{�4�B�I��s�V������ �5��[y|";
�C2O��.?�ȝ�G��p�9��Έ�5-�q
3�Q�NY5W�@}��Mz�ћ�;�A�	�E���H�
�M 