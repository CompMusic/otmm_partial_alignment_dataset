BZh91AY&SY݅� f߀Px���g������`	�{q���I@ ArfT�JT$P�	1�Dɚ����⁣#L��4 �J��щ�& �104d���`F�b0L�`��4�� b�  OPѓ �`A��2`�D�4	���OI���P��Q�z��c���H�I�E� �~dWrbR�P j!�����
D�����)�����t�JQլ���h�^fff]���fffffffff.fffVa��m�1�,��]���`مk:#{ڒ!��D[�M[U��ۊ��X�5ѕz�h~:`�)2�7g1���̫2da@w=�}F٫y�|(22d�a}2��4�Z:�gFF��B��+����e^,nѳ�[����7�(� VJV�	.k��Ei�R����OQ�ը�N�+"F�0��"�"�Z�
�$�" +X 4���վ�?,�Ief�&v;.�����{�j3��WDd�	8��2�vA�]734U�b�W����s310�6L5X>���6s�z]V8ʋ�?�l�uj��8�J���㵑�E��	�:��7%�D�$	|���QuVl�:l�i�j�ZƎ�l@۝wx�E)��v�K%[D'(U��
�p,�A{�c)l݅@�-
���SY��;INKn]]i+p9�l��T]ε����e�]_W�'Rp�r���h�d2��A�p��	��a����x�&(ç-[�NU�RI\t]��	��W��&�E��xu1?�0�^�-B����B�Cc��Uj�v+U�-wM�y�C&�6�Ķ�;�>^cތ��J�5�dd<0uBA���05m�q�,Su�������Z��Xj՜gvw"
A-5D3��� q0�\��k�Z.(�@�F�����w�J�3a��s��U͐ܖ91gx�����7��b0n�������T!�J�,���_�2��.�op4_���4'���3�/J�S�T�T���)�X�d�Cj�8>I���ă��� t���K�d'Q�(�{��pG������j�a�������B�sZl�����s� ������b���_&J�D���knh�fV����U�:���f��<�^�l��ِ��'�DQ^�m����͚�/Z!��R�T
R ]�����`�*���IL�vʒn�pʑY!rQ@�"�.��J�ZT8��� Z*�B�87ze')7��mX�h%)v�Q�"�\�"��Gw!��^-]z������-M 6 6Z�ь���s����Y�&�"��C����3�S�˂���D�/ns�/���0�G�* ���ݮ�����"� x,Y��y�����ͥ��`iK� #[  n��笎�۔ù:��Џ� �ּ�l:q �W�{��� �ٺG�1��ˮD�D�B���o&�	A����x�^6{Ĝȭ,�V�y�j����C���k��U�����I���U�`�*�� �4�)Jj�Q��Ӈ����]��8Lɞ̣a�GN��0 ��(r�jE}�sMzu��Y�P��t��!�H,�ea` ���T�Օ��x�nZ  �@:���|m
r!�9DՑ�+��B��bE:!�6���t^RqDy�v�+�wW:ܷ�!���5���N$y��]{�ՃH@ S����/� �k���J؈���(�G ���rVf4`����4 a2520mK	I�A�����q�Q�u��0p�����B��x!ܕ�jL�2�ANʢ�4�&u;
 &�F�Y�wZ���9$��ĄX�a�XvZ��X��9�a��ݠ|-����5��T�B .�9&1o|�� 9�gô��,�;��/ʬQF�ni3����i��֦�1�V�7�h�-�BY��5�S�MF*� w�D�'��H7��ȴ$�zW0 ���l��R�\h��������΂D6��@.ꊳ,%� �(΀	:�9O6��nT���c_Î;cٌ�}L.8Q�VG�.�p� %��