BZh91AY&SY�r� I߀Py��g������`�,xڀ  �ܒɉ�BBH�4�A4ɓ�df��@�2� H�6��� #  �� ���&L�20�&�db``��"���M�4�   hsbh0�2d��`�i���!�D�'����OQ�i2   ��ed{u�%�D��bӦ�-�'O��_��(D`��.� �r	�B�d�T;��q\i5p]�1կeTU�d�痙���wwSvs3.����3/P\����p���>���^�O]��J߆Qv�iql��`[L��#M���"Q8��9�ڡ[%�#-k:���W�}6?k��?<7ўA�}�Rcf���2+wf�[[�$fV�eޅ�ݢ�2Y�L^K��[K�百x�@�l�b	����ydr.5եTx�#�42�[ĸa<�	���mdL�Vj��j���00�f��椉;���C�@�]U�ʹVW#��%����o0ق�V���2P KT\�,����UHV�wARA����{)��+�g^�)���u3��)�08��k��H	�RZY(������� r�g)@YP�x@�BR�$&{,�
��0�z(�����M=Xq�#���e�Yq�3nI�+!�.Ǒ#�ݦ�snC	"��hɪ��wY��#��*�,�W����49�km���n;��(�h�4�S���ԪN���I���w��z\X;��lVL��i5EB�⏽>�����v�-�r{3=#Ȏfs���㉘�f�#���W����R�u���W�a�Hz�	�5T1��8R�*�LOSЀ����`�47'�	uRȳ/O��D:���Ű����g.bO"�q��	`�q��Pj�W�nR-(K�q�d�>+��*�5��R#p��~�b��FCGYˬ��uƆb���h��)��Q�
��{#���A���7�J/]�@�k�6
�Ha�)�QD���C�N
`��cԛ�0�V��q��ĸfKɜ����RC�g9��|�j���EN��Wb�4�o�6�C2,�;��S�DQ^5iA*�`��>�m�dtX��_ UbaĉȒI���*$Ȣ*#B��*IB!S�<c$�֕E��q��L󵒲ȕ���B�B��R�;K���Eګ�Z� ��[48�a2��G��ߋ"�!��od$���棤��k��o�"��H�Q��R������Į�������i�7OLO�U�["{��:�]J\e����:�;x�8���X�ESdT�Wk@%�G<�[�e`��'AO~tG[��� �R�B�)m���%2��4(��#ZM�Mq�6����ʊ�����W���uƢ3�lã�����ka�sǀIZ;"r���Dj�h�UPA@!�TeK�(d��7�(�8�����4D�#ƈѤ|f����ǵ�~��v��՗n���jD7(�B��L�3�}	3�� �7�\� ɭ��V�ٍ�[�g5�}5�gm�t$e3Ȱ�����j���3��D�t!XHL5��D����=�Z+��3�HZvO�'WY��D����Q�+��@Ў�A�`���c#M&��k�X@�n�{�b�:l��+E�r�V�*暡K�®f���.Y�B� ��r/B|�R;��Z!'`���nn���#��be��On�y��|��)���� A������6P�)|�0r���2�m�/	3&�p��A�6��5���50g4U�E��W��%��^l�Ѕ8,��dZ���e��r�A ���;�#\ɲ��,8H
�$�g���G���S�+��QXi4i�(��z:�@�paxg�B?x�!�N�Q�	�"���ܑN$)��