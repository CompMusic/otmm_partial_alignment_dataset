BZh91AY&SY�ԩ �_�Px���g������`
���>�S��  ;�}�^n�m�wiP�Dd$ؚi����i�ih�4Ѡ5=Q)�!� � `F���F5 ���h�4��L��P��
��4�@  h L��IM�D=OS!�M=C@  4 	�b$�!�d�   �s1A#�(̂��B
H2�|��I$<��H~�� �p$!�zX|\�$A�	�m�����4�^��'�y3323ff,̬�|�����332��UUe��ä�>���r=�\>WY�u����i��]r�\�2Ă��[K�!;�J�����M����$�{��Q.���+(���˶�����v����rm?6AB�a��'���a�F$�*g���V�T)-�j-�	tPR�LʻZ,r�,Jq󙣫~�����{7��$��LE+�7��+����)�Y%�ԩ=V\d���3e��m���p�Nc�TqSkd�P��T�	 dɆk�v�`�焲,�t�1,���{x���[����J��W�NJ3��eW)�+f��Kj�j�0[[���rȑ��!�pj�)m��6&�¡|bܞ��݆f�2t:0��������a�P�]����'�!��>Y���Q�90� ���r�hy�u�0��A`�(p65r[�8z�^ķ9�7������5=�ku�L���)a�QD�w����������=��	���̿"�Ld�=䫖��ѣ%� �y �0��$r�4��	4�,CK�D��Ŗ�,�e��9,�J	�Þ���Ȋ��Y�]�O8����}ŵ/�F8�7|
N)��T���/W���T���!�� ���{�`���t4�<T�r H\���]ք��̓}|�4�.<lk2\U�k����4��W��E|Ar{$=:mnˇ;B�d>0(Dm��z�&���/E�5����������L���8f���"�.e5G&h8D&�B�^�`a?7��Dq��1��"�t��ȧ��Ζ)A'�Pg��_��vH, ^���fW"�4�B���"n]�������`�1B��N?u�E��-f�mi�azs��=��y>6��s��y�we[��7h�͙�u�.���C�wO��虄��(��"u3`�8~�Y��I�b]}c�q�����p���/GϞ�	^}ȶHS��h���\�څYȗ2�@ۅE�&uE�;:��֚��Ǡ��	�q@�Z������é��S0[��š�m��I���v���Rxޭ����$}D���@�f�<����R�T
1$(:�j��H�����TSUPb���<�Q�<�!L���i��TYYH�ʨ�zhi@8�w!9K*���`-JuŖ]B�B�cAXr����<\h�=l4!�;>���
E6΀$�ЦkH�Q"�8��dL��;&J�e�W�1��E
8��K!��vI�*�=�!�۸/Zr�RP�ե~���d���_޹�"�Ua��T? �e���s^S|Ҫl$.$e����1�O.`+Rn"H&��+O=�˒�_%f��c*�KOA���A�{V<u�X4ؤ�͒uݽ�^��пS��5q<�bQ��g��n���<�{?f��1`C��ꠈ�,X,b�+�h���((�b�`*L��	Nx8���s��!�z�\K�-�P�RL
2�M�V�~�u��(������6h�q �����$���m�KK7:y�,�a��$�ptY���_z�:x�sAd��9-%	�wfk��j�Z�!I���S�Z��t�@�`��Hj�m�o0�{'�n��4��9�^X�D��$��]@B_�,�%(K������EC)cEd%���4�h��hF��81�����Pù(2x��C��ce�T�$¥��s2bt�Ψ׭�9�-=7�D�FSl�&��V$��Iw�H�R=���þ�ɜ2�jA�[��c/^q����<�g��r�J�N�H���*�Pv^�M��u]pl��d�6�sI���r{8n�E�^��E�1�F��
��Yh��*QOz�v� �]�,��P�p`Z�.�&����)#UdL,K4�Q#N_׌��I�6���}jfA�`�[�F�nb�I�FĒ	w@o����ܩk+`ƾq�3�:����M.�ŋo�]��B@v3R�