BZh91AY&SYk�� �_�Px��g������`{suٸ� A���m�$B4h5&�=I�4G�������@�        昙2h�`��` ���M$D��24hz�  �i��&�&	��0`��$H"h�#ڏ)�H�� �K��Oݭ!�@�!@��!���$��V�>`?}	�@���a!P�2��l�nQ�7�p�<�9�s��9�fef.fe����ށ����.�=��+�p�Ufmy�gp�A%CJ��X�0��;:���t��S+���d���Y�[lϬ�(//d��c�tH�-+@�;b�jw^�WY����q}�5;���RHW
�	����+��곫W�g�9J�K��+Χ[�V삥�V�*+Uj	)Lʶ�CM1��]�7.[`68�Z��L��y��9�1��k3�imӬ�)�;��e7f�[Mͺ�-P"�Uf�����H�IsL���Ս� ��.��a^͇Vq�z~@0O,�C�6���)�@Σx�h�KP����q�df3�Vm
t��Ѵ�N��M�����I�N����rÁ
���tU��hn-R�!�I�4/1�XP1BT�8Bhu<:^��|՗C$�����y�hJ�lĠH��|��[[QN��9�}�_yˈ���届N���-J�"p4OZ�$M)���p!��1�m��C������e�_脡㥉q��!�<��'9#i�H�G�b+\�@��m�k�*Ն���Re�W��Y��h�qF�VG��Q]�r��Kf�&�VC�+7��A���'�ؖMl5�ӷ6N��$@r!�_X���mex��g�^'[�-�V�X�T�
�Hb+���H��L�m+���׀Tg��q� Tg	����g�x�E着$&x=��yLcu��a�$�wǔ�_�.RPQb,z b�Ѷ�cK*���j((�*Z���;iPގ0��`#��q�x�Y9�c�
U�)4Q�h������ 3f*e7�k�_�QȪ����w5��t����J��D���]؞}�5M�WC�'���*g�}�OMP���E����5O�����H/KԄ�׶#� 7�e8=KM��5&�I~��h$c�zby� ���	���=�>���bpn�4J1D̃bP^�[y�4�(3�|��JX��vb�Iԋl�r�A#!�G;+\��RG���ξ�^V�,�X�d-����*9�qVX��'�P�V#��\V2Q�$'L�N��`�5fL�*t��u��]z�b���`����#
��`��}i�Ã!"��-Ԍ��jѱDn�lIR����GyH���#^�寁A��"%�3a�t\���ˮkh$Z�	6b��� o��5�]s�2ݵit�w��L�:H�#��r���-NIM�`���(Q�dX��t�a!��}D�"�ν�5�	;Ǉ�`n{^���npz�ڢu�!ܓ����2�O�b�t�5;JC&էG{�h'��i�;���̀N�����L;�_&q�e҃��!�0ë�~p��H�5=�ء	��oLb�v�k��@H���SU֝8��
��V��*��a �$����%�U�9�|��ق�_c�����*Tb����H�<]�j�0j����@8�YD�q�$��)rD���bE��~�&�����;�-4+�`Hۺ��f��Б�� l��LK���kR��[`ƾ�3��d��/��r�w�.�p� �ٔ