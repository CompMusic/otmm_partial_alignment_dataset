BZh91AY&SY�.@� 
߀Px���g������`	_,{�����
�_|�ͨ[����	$L�ML�ѐh��=C	�'�i�A��4�*P       jjz&�Dhd� i��i� FF�%=$ RM�z�@  ɠ @6�=#MS5��4�@  ���� �~��l�Q��4��� 44b=54� >���$ ��E�  ���Y6&��x$��R{��L�pg���@E�
_���ãf�B0�vͰ��)fffffdDDFffffVb�fffVb�h�n�B����@�ݤ���e[�&;�4����KP�j ���N�)*�DL+Qf�/�g��ǘb�e$&K�c�l��vV�*T%��'�֦k����%�4�p��$�b_l�fn�Z ��j*ؐRmЁ[^�#8$��P*��etL�6#�eLݟ}t̔�эn��i�qP�	��H���N�"�9���@0�&k�4�vLO1c�z����;��[�X�~}�^�K�&/L^2U�wŮ�&�-dĨު?pM�� ��y�G�瀊�D���4/�^�4��!��j���� M�U{]\��QI�nyߍP��E!���5��g(rBfβ�0˨D��z\��V	�u�Y#��eJ�M�k6�܌��N�w�F�s�	@���YQJ�H��pb�ekJ�Lg�w�m��P#T�-a�=f�t���J�\��|��@b�!��HTb�9T֩p��z��K1�"���ٕ�����vB��ū���x+�bȒ���1u
�:P� �T
t�l��O�KwĊ�ɜ`��\;���R#�D�+lH��qs�����Y]�J�E@̆np��!M��F��VrzTp$�+����>
Khdq�����b���	�kb�łդLqpQ�i�u�2��U�s!Ux��:�9.b�`�ε���xf�%��8fj,@�g��"T5��L#�!Ӏ�'�'��F�pEFo Uz�3W�r���l��í��2.�R���Ec�N,��Q�C3�%Ya�t���]G3����]cT�R������Zbm�釐���+bZ��eHR]9<Z�����H��ƶ�4H�G_�h��=]�[7�vvq��{�=UE{UU������^tB5�R�P(�$⃤l�
i�e�F��f��oFؔj�0�K��jbX�Р��b"4Ҋ4��Ugy�j�֍��B�K4��DE� !����k��E^F�.k/*��`�e�v@��6�đ��{�xe}J�nӢ/�F��`4	~b]������L]	�/d�r�u�MZb �ޛ�G5}{���$�2^��j\�IN���[��Y`l�V��e|\�	y%�B����m+�Z%��7V㊙_ܦ���0�U4�̇�2(��O�t�L���h]|��yQ�$�<h��A%I�[�����:��CTW��Z�j�JQT7���e �r�N:fɲNq=�����i�b�J���Bi%���<�&Y�o�l�v��76�G��\�`I~�B8��t/��)w�Ɖ�	)j�C����dt���鴍
���bi��"�N�i9,�]9H�0�3�;�l%��K�32L5G&ze݄}�p`����ƀ�����+d�˴�K�Z� Ȳ�3��dV�
H�0Kq�U�3��	+L��L��+L(<� c	�m�,��V�ce�$����!He���P*HC����BI�k���p'���׉4��# I���L����T�A���5XF��ѽ��������^D�rR��0��k���KhL	*���
�ۀ��`���*(�m�&k�@3���{i4�u=kS�M��E�7�`����THԧLȧ;@"$%���B��(^����B�t�� &S����TӜ_͆�C��N�������@kpEF�
����h�uɪ�<GaƩs/�ƺ�j�i!hIK ��]��BB��