BZh91AY&SYZSѬ ;_�Px��g������`��� �{�N�U�7�IOD��?M)�	2x��1����4� ���H�    h4 �I�j`&	�CCL�4�!��@�	OI��x��H4z���� ��49�&L�0�&&��!�0# �!4)��<�m#ҏP dd�M=K&�U.�H!4P1���2 ��=�M���%�!C�O����`.��
� I$T�������y<����yw33+0�f6]�����ff^�v�ef�<aý�t^aY����+�<��F$�z�H:(��K���WwhV���j���E��<��ɐ���1���ym�н�d�p�Sd�'Y��9pȈX5"�{���.�����W0R�k�/�g�������M���qE$�%l�]e���J��Y�p��c7���}>�#%��>~P����V���`��E1f*��H���pŘ�.d6:Ū(�V捺����s�d�$y��z�xpVJu��2�b��
�űP9��W8�
�"����{! u
�J��n=E�F��[鱒&*�zeQ�����K�tB�҇-`O(r���j�ٷ�dǈƮ+Z2�	�_�UE�4��
I��Ά�2���#�a�v����a������sck�)�H�8,�6�PW���
��;��N#o/�q8�Pf*�P�(KpAUY���� Ȝ�U�(��fݑ�d��k��6��\c%��q�͸*���K���qS�Z�(Q.��9���]P�+%>�R�TVN�2�D�B�e��������s88 8�c�:@������/V�k���Ed��f&
S>���ヵp�8�gz��g��R��V<(��L���������u�t�M��c�7��9V�+�v��+�UX4�8�g�CM^���*�R%3ڸ|({����(���Q*m��o���芊��!AiR1���r�Z̄��Q�E�f��$sp�f!�!�B��ZMx4Pak_j; -j��Ty��ś�XMH�X��%�b5XA�(i���`��g��)�8vK�Q'55�5l�W���U�/;�m�'cOJ��ލV���a�\��6l��������h�u��&I�K�D���g�@���*�x����Yi� ���2g�$q��m/)�)��"jQM���߲R�+�n"OEI[mת�!���ʌ%$]�=�r�:�M�ɸ�PZ�E�=ċJ���G��N���*��'ǔ�P�����J���!-EU���MjV�"��pA���L:�
�8�L���D�x�]7�?5�	(�����qC\lMtr4ׅ�{q�Ɠ���:��T���
LUPq�fwK����Mn���H"�ث� ��L^l���mt��R	t�@*�#��\�h۴�ƒ$P֛����)	�K�-ТY24�2/$_�@�X�!h=U�AE�<��vh,x00� R��+��5[�֓���S��Z��E�f���C��;-����M|D�߳)�T�����ߘ:�D7;P�4D<�=�=d�H��D*wN�	��n��{�!�A���݅�_�݂�� ���J�-+���� \n�9�������-�~��!2���J22��� ��a���,���%��� �טY�����D�`�Q(��uR3��6�&��E(�&d�\�d!��,زĹ!MHD��@u���>��J��5�ơ�c�HY���@�����"�(H-)�� 