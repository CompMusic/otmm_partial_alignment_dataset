BZh91AY&SY�U"
 {߀Px��g������P��Ɖͮ95��w	%4)���)��A���hh h�&���4'� ��� �d���O)➐4�@ ���昙2h�`��` ���H��T�=S����z���� z�(���$����" W̅��16�@�s���:hp�^fM��� .kvskӖ��V���9�inI��ʶ�|muq6�����P���:	�%CS gX�0c\�jO
QTo�Yd� ���^�T��)]��`�c��B�`-���<�-L�fw8$ލ�.��A����
��1�s_q'-B�U�d2�Ú]8����������g�]��\XU��!��i|�����jWJ������66�m��73S�o!����EaV���fGC�륕V�축�e�0�kƫV�V����Q��c�he�_����fG򈾩��՘�4�v�W��Bě�Z՞�F�R��'{�av�_�q��s뢹�*�Er����ƍ������Ό�c �D�#V�_�s&�3�aKQL^��-c�[����j�@˻�8������M%lh/A�p���Q���!��Ή}V�P	L,��(w�gm"� �F�����Z���70�x┉<h*:�qc2e)��L.G礼�ag�Իܺ�.%^���|
n�X�P��3�D�ue��K��Np��	&#�)���#:��vr(��5(���HO���U�g���6�X�p�N�r�`��J��L�p�9�k] �g��瓡���X�+(d�G��x�de���.7$�G@}̔��R(:W����0��?-@�/`R1��	.�����������¢V�V3�Y䉨���ՄVrs�Lc�9�A��򈁃g>|����=p��.�N=���� Y����hxd��~���4 z�������7.+-(2�-��tI�v�e7�׮2�!��4��b�V4/~j�L�,U'����\��z�a�����$7c�e���B�+�!T�W�E����a6�� �hR�Ҫ�ܻ
#nD���)�:�0˃=6?T��X+/�w$S�	�R �