BZh91AY&SYn�: W߀Py��g������P���;��z������MqxID4ɵO&B=@P4A� $��45i4����i� CM4��j&�OQ�i�P4 h �)L���Q�� �M ��$��L555<�T�)暧�zjhhCA��Si���P&��Q����I�F?�2A�ń����݀�DQ<e�1	�Te���gd�znaE�$�+M&(����%��#�i����!�	բɁ}°(1)݃�H0��j#��M4垹ڵ�Ȁ�̅=M���� ��b���,1J=b[���y/e������b�q��N���<8���,T7�`��s�iN��R�%�S���K��5up�tE���D{m]Z�=0��&m�ѲU	�C��+��!�*����d	p-+��DWL��"��(����\�q^:l�������ۣC��w��vHBBHp�$��x�����2|��X�0��Y*#q�◍�RN��(�3�Ӎ��%DL��R��ji1�Q��F�^j�\�45���W2+"�D74��ӵ�ڬ-�%�X�zhovC"�	�.� ��@z�<��UA`<{PԠ�j��#I�d�m�F��]j��(�S@K���+*���P���R���`��cy��1V��f$��Ե�x^ue_��-yP,-M�ͭL�F'FKБAI}����alvAj5�0|�lY���nA呼Q�[u�D[��(TTc�KI����(��s����M$�4I$�	bSb�vA��0�x��LE����ff��^1%m47{���.���g�έ^�!�bPQ-L� �X�����ܙe�$H��n���*II�m��W^ƨ}���5�d���m�mgq	�#IR+�VB�dp�ұ�Ѓ0�,��+��X ͘m&�;3^�`Gë+�& �_!V^hJs!�0M�RZR�Eܓ�k|�	���N�δ�ivŕ���U�)m�b�v4X.����`-�DԶ%T2{":n,�,��i�(_�@�`���s��p��+rJ�c��o8��?y���!��x�#�r�]�C5��~���܊ �[/�q@_��pkOj���(���ޯxQ�V*h���HUX�P��u�2e�������
{���M��`�c�!��[���P	Pl��̒Ж+d�khZ�Y�bL"�y:���$��HtB��SI[��������G ZB�*���p`]����_���r+��E���B?��Rhw�H ,߉�#�W���)��vY�