BZh91AY&SY���� ;߀Py���g������`	�z�;ױ�xl��hdi�HI�����zyS���6�G��#4��CSA��J�P=@   22 i�	�)       �H�z���4�d i�4!�`�1 �&	�!��L��JSК1S�țI�b��@i���dd=L�@oJ(p�`��Y�����3lT��H�0�s��Ք@Ā���!}(Ǐ+��7�캪}_[�עI$�I$����I$�H$�I����2��E�!}��xO����ш�ws&	�r-�����tB�����2t�<3�.�I�j�o:Ѣ�m]f�#�q]����-��54C#�d_G�����:i3zf��W-�b��������6/�x�t�)�Ȫ�f�5��q���w4Ջ�vn]&)�yh���(@!��6���(��9Ӕ��J�)T<����[A$ɐ�m�|������U��NZ�Nb!�8A��6�ic�c�ә�Z��[w&���m��YM7.�r���_�sN���u���S�8⥢�f�j�RjnD5[<tc������Mpb,�[w�����l6'M[�4��0��$�Y;hYQD��,L\8�YgX�����}��'d�^�0Pt��n�+gh$�� �0ZHD��8-��}��1�N�����=�8zQg�q�9�) i�g^��(�xn�VL����j��j�Rz����vl�-j����<�]w�F�m��D�`YS�z��[�,l�Q���gb� ��ࣗ�+v��`=  ��f��нƛ�!�7s,�3�����uJ�r ��~�g�*l�.)[��ȨqɍP&p�"�b��2Q�^rZ`�M	ӆ����Rӫ��y�8��sh·%���\*1ppj�^�>%�7721h,Yv�v�ԼaOU.-�R��\*����n��hq�Ҫ��C�H��7�C\!��P(r�"��VŦ���[�;�Y��q`��\[S�6�)�sh�E����hf���Ӥu�k���;����ԅ4�_�x��0��w��
w.:Hm�]Hٷ�nܨ03%�6z�e����Y��,�U.7���\
a�0s�M�^��⳷"@xƔ�ϓ�y�w�@�A �vUUJS��v@�N���f�f�I.f�|�>d�m
�H�JT�)�*��P�B�B�]��
 ��1N68b݁�	���c"ά)��`����ŤV��'D�Vt���':�u�hChs,2q ̐���V�0�~���V�[іH����Ɲ��}�d��N2z�b{�}l��WR{ZQ<{�*��Χn��,����bc��Y��+x��4D?�+��C��8����$�r��q��Ff0�U�`�_A���KC�y&Y�M��_�$�l߼}�ܿ�/�G�f[!z�:�u���#�h�#�אX�BB�V	���a{���b�='R�9�J��ۭr-`�t�ۺ�
g'���c ȒH��FE� ��k&І�� ��rP�B֥���%���LB�W�F(��b�m\�9�,r�;D�6dzu���&���7y�pd
��(��>���>�)L;��0��V��bw�N�S�v�S�m�f���j��EvN]��֡i�?^�ġZfYE�(�`iԏ¯�ެ�/�ŴW��������X7e��'�;�{Rm�VJ�c\Q�W^�W�w>D��)��֑5�,�y� W�pva���]e�sEs�l�#¦~뒅y`(z�i�4i;}^��78
4���T$|h�b8%�Ǒ!�jp�1l��Ct�.ahk;ś9���m,��͠� ��z��p-�ڻ��ZQ�B�d;��F�hް�{�v�J�=F����'P'�F��6���V����/ۗ l;���{)�8��З�˖=:��VP����gMI�������i
�Ƞۉ��,T���uA%5�ĺD]Ǖ��`ƲA ��±ЪU�%�I�l�I��-�C��M���3���
�1@�O���1�+���ȭM���h��`]�1��x��_�	-BR!R��.�p�!����