BZh91AY&SY�[ �߀Px���g������`���_^��!�j��=����ƥ� =��M4d��Ѝ  SA����i�0��4��CLF��IM5=O(Ʉ hM41����P=@4i�   @Ih��h�h �  $	��蚞��4�=L��4􍩄�:+j]�j�:��"�j ��I���*��	H}l��� ����� Mo�b��~�1�s|��G1M4��������՛������5UUo�M̺��[#�K�I�<�\��"1�Ɨ�5c+v1d��;cgYAb���V�L�I�#�bq�6dv]��z�	f���"�BZ2|�cL��fOa2r���Q7��$��B��H�Lüh-F����r� )�j�3M�k�h*y=��d.�����N�C���Jp�%a�z�4Һ�SN�A��,X��M1���u�Pe�K5��]=W`���è8u�ځ�7�d]^ K�:�0�;�cS�R�Kg"���o�0;+
�K#&\z��G�H�����V�I�+ҡ�4 ��&����A YG(A�pxE3E��e�J��0v}��3m�`-�Yԫ�-u��Au��]FZ�s{���Pʈ)6�s �� %ĭ+��E���1�p�Dd�]FY�Dˑ�@v\��@�u�I�It�ؐ/e��|���U����dSDl��5�iQF����*�(E�>Ԡ3V�]$�Òj"U����i34��:����me�c�Aa���vQ�D(җ,���ڢYA�M���Er^�[�}p�'c+dr�&�[B1c .�n�1}���5ZȴQ3CJ��tn�����nHui2�+��xz@N�1	�r�������%b�e����|tpcӚX�#t�5���a��1{V5z�����D���99Β`��Wނ�Zt��'�4B���oo�8�nmMh˲��7��LB���M�^���� �
mE�Bm�dH4��^��@c �`���wܫ��wy����ۻV�iw���Zj��ީ����j�]&�mQ��4�:g5������Ew*�	�����C{�+���	1V��j;�a�-
U�e��5GT�lJ,�j��T���M06�%Ҙ
cmt� ZB��%��f�a,����"�e46lf�/<�]��kV&�كW��G��:�}&�:�Ԧc��;~�>�+�Z�'��ػ7����⭐�Rg�� �MM���=J%@�z��u�V�I�y4�xJK��ԙ���e$H7����p�����M��H/�'�@�j�2�����U�������#����#$A�h1Awr\�h%>{/o��)|��$��J����,�:����m�-h{�>|#7���x��h*�AdE�AH�MJ��B�8����MU�d��~�E�$wq41S&����5z�Ms�T��hR���KF��t�~os�P# ��Ē7S�(;kն��Q. H�]��F��WlQeē'��+���o�n�	�v��)U[	ș��!�m)�^��K V�$ǘ�\9i��<4UU�m���!=尪���/F��&ʒR��1CZb
m���x����5!-�YL�[c#&Բʀ�f�3��]�jHE���B���*L�˦�3�1����h��9(	2F�5�8'��f-�� ���C*Qa�ꯍ!�̽�V,n3B�ǧ����<t;��^��J�
���+��^^0�`%C��^_��i��E��ʊ6�r$�q 
.�۶+����a]2�<�hsX�ł�i�;�	W}�;���݋�2� ��y�x.]����	
����ѳ�����%��AxG:����Xq��R���	m�&�)�366�ゥ��F5��g�g4-��=����w$S�	 �0��